// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_044
`define RVX_GDEF_044

`define RVX_GDEF_171 15
`define RVX_GDEF_213 8
`define RVX_GDEF_341 3
`define RVX_GDEF_321 5
`define RVX_GDEF_015 3
`define RVX_GDEF_051 0
`define RVX_GDEF_142 (32'h 0)
`define RVX_GDEF_127 1
`define RVX_GDEF_205 (32'h 1000)
`define RVX_GDEF_025 2
`define RVX_GDEF_347 (32'h 2000)
`define RVX_GDEF_359 3
`define RVX_GDEF_426 (32'h 3000)
`define RVX_GDEF_065 4
`define RVX_GDEF_262 (32'h 4000)

`define RVX_GDEF_353 12
`define RVX_GDEF_391 3

`define RVX_GDEF_246 12
`define RVX_GDEF_064 3

`define RVX_GDEF_350 12
`define RVX_GDEF_147 3

`define RVX_GDEF_374 5
`define RVX_GDEF_283 3
`define RVX_GDEF_121 (32'h 0)
`define RVX_GDEF_111 (32'h 8)
`define RVX_GDEF_259 (32'h 10)

`define RVX_GDEF_257 (`RVX_GDEF_426+`RVX_GDEF_121)
`define RVX_GDEF_138 (`RVX_GDEF_426+`RVX_GDEF_111)
`define RVX_GDEF_033 (`RVX_GDEF_426+`RVX_GDEF_259)

`define RVX_GDEF_220 4
`define RVX_GDEF_129 3

`define RVX_GDEF_226 8
`define RVX_GDEF_242 0

`define RVX_GDEF_207 11

`define RVX_GDEF_084 11

`endif