`default_nettype wire
`include "timescale.vh"
module IntSyncCrossingSource_4(
  input   auto_in_0,
  output  auto_out_sync_0
);
  assign auto_out_sync_0 = auto_in_0;
endmodule