`default_nettype wire
`include "timescale.vh"
module Rocket(
  input         clock,
  input         reset,
  input         io_hartid,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  output        io_imem_might_request,
  output        io_imem_req_valid,
  output [31:0] io_imem_req_bits_pc,
  output        io_imem_req_bits_speculative,
  output        io_imem_sfence_valid,
  output        io_imem_sfence_bits_rs1,
  output        io_imem_sfence_bits_rs2,
  output [31:0] io_imem_sfence_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input         io_imem_resp_bits_btb_taken,
  input         io_imem_resp_bits_btb_bridx,
  input  [4:0]  io_imem_resp_bits_btb_entry,
  input  [7:0]  io_imem_resp_bits_btb_bht_history,
  input  [31:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data,
  input         io_imem_resp_bits_xcpt_pf_inst,
  input         io_imem_resp_bits_xcpt_ae_inst,
  input         io_imem_resp_bits_replay,
  output        io_imem_btb_update_valid,
  output [4:0]  io_imem_btb_update_bits_prediction_entry,
  output [31:0] io_imem_btb_update_bits_pc,
  output        io_imem_btb_update_bits_isValid,
  output [31:0] io_imem_btb_update_bits_br_pc,
  output [1:0]  io_imem_btb_update_bits_cfiType,
  output        io_imem_bht_update_valid,
  output [7:0]  io_imem_bht_update_bits_prediction_history,
  output [31:0] io_imem_bht_update_bits_pc,
  output        io_imem_bht_update_bits_branch,
  output        io_imem_bht_update_bits_taken,
  output        io_imem_bht_update_bits_mispredict,
  output        io_imem_flush_icache,
  output        io_imem_progress,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [6:0]  io_dmem_req_bits_tag,
  output [4:0]  io_dmem_req_bits_cmd,
  output [1:0]  io_dmem_req_bits_size,
  output        io_dmem_req_bits_signed,
  output [1:0]  io_dmem_req_bits_dprv,
  output        io_dmem_req_bits_dv,
  output        io_dmem_s1_kill,
  output [31:0] io_dmem_s1_data_data,
  input         io_dmem_s2_nack,
  input         io_dmem_resp_valid,
  input  [6:0]  io_dmem_resp_bits_tag,
  input  [31:0] io_dmem_resp_bits_data,
  input         io_dmem_resp_bits_replay,
  input         io_dmem_resp_bits_has_data,
  input  [31:0] io_dmem_resp_bits_data_word_bypass,
  input         io_dmem_replay_next,
  input         io_dmem_s2_xcpt_ma_ld,
  input         io_dmem_s2_xcpt_ma_st,
  input         io_dmem_s2_xcpt_pf_ld,
  input         io_dmem_s2_xcpt_pf_st,
  input         io_dmem_s2_xcpt_ae_ld,
  input         io_dmem_s2_xcpt_ae_st,
  input         io_dmem_ordered,
  input         io_dmem_perf_release,
  input         io_dmem_perf_grant,
  output        io_ptw_ptbr_mode,
  output [21:0] io_ptw_ptbr_ppn,
  output        io_ptw_sfence_valid,
  output        io_ptw_sfence_bits_rs1,
  output        io_ptw_status_debug,
  output [1:0]  io_ptw_status_prv,
  output        io_ptw_status_mxr,
  output        io_ptw_status_sum,
  output        io_ptw_pmp_0_cfg_l,
  output [1:0]  io_ptw_pmp_0_cfg_a,
  output        io_ptw_pmp_0_cfg_x,
  output        io_ptw_pmp_0_cfg_w,
  output        io_ptw_pmp_0_cfg_r,
  output [29:0] io_ptw_pmp_0_addr,
  output [31:0] io_ptw_pmp_0_mask,
  output        io_ptw_pmp_1_cfg_l,
  output [1:0]  io_ptw_pmp_1_cfg_a,
  output        io_ptw_pmp_1_cfg_x,
  output        io_ptw_pmp_1_cfg_w,
  output        io_ptw_pmp_1_cfg_r,
  output [29:0] io_ptw_pmp_1_addr,
  output [31:0] io_ptw_pmp_1_mask,
  output        io_ptw_pmp_2_cfg_l,
  output [1:0]  io_ptw_pmp_2_cfg_a,
  output        io_ptw_pmp_2_cfg_x,
  output        io_ptw_pmp_2_cfg_w,
  output        io_ptw_pmp_2_cfg_r,
  output [29:0] io_ptw_pmp_2_addr,
  output [31:0] io_ptw_pmp_2_mask,
  output        io_ptw_pmp_3_cfg_l,
  output [1:0]  io_ptw_pmp_3_cfg_a,
  output        io_ptw_pmp_3_cfg_x,
  output        io_ptw_pmp_3_cfg_w,
  output        io_ptw_pmp_3_cfg_r,
  output [29:0] io_ptw_pmp_3_addr,
  output [31:0] io_ptw_pmp_3_mask,
  output        io_ptw_pmp_4_cfg_l,
  output [1:0]  io_ptw_pmp_4_cfg_a,
  output        io_ptw_pmp_4_cfg_x,
  output        io_ptw_pmp_4_cfg_w,
  output        io_ptw_pmp_4_cfg_r,
  output [29:0] io_ptw_pmp_4_addr,
  output [31:0] io_ptw_pmp_4_mask,
  output        io_ptw_pmp_5_cfg_l,
  output [1:0]  io_ptw_pmp_5_cfg_a,
  output        io_ptw_pmp_5_cfg_x,
  output        io_ptw_pmp_5_cfg_w,
  output        io_ptw_pmp_5_cfg_r,
  output [29:0] io_ptw_pmp_5_addr,
  output [31:0] io_ptw_pmp_5_mask,
  output        io_ptw_pmp_6_cfg_l,
  output [1:0]  io_ptw_pmp_6_cfg_a,
  output        io_ptw_pmp_6_cfg_x,
  output        io_ptw_pmp_6_cfg_w,
  output        io_ptw_pmp_6_cfg_r,
  output [29:0] io_ptw_pmp_6_addr,
  output [31:0] io_ptw_pmp_6_mask,
  output        io_ptw_pmp_7_cfg_l,
  output [1:0]  io_ptw_pmp_7_cfg_a,
  output        io_ptw_pmp_7_cfg_x,
  output        io_ptw_pmp_7_cfg_w,
  output        io_ptw_pmp_7_cfg_r,
  output [29:0] io_ptw_pmp_7_addr,
  output [31:0] io_ptw_pmp_7_mask,
  output [31:0] io_ptw_customCSRs_csrs_0_value,
  output [31:0] io_fpu_inst,
  output [31:0] io_fpu_fromint_data,
  output [2:0]  io_fpu_fcsr_rm,
  input         io_fpu_fcsr_flags_valid,
  input  [4:0]  io_fpu_fcsr_flags_bits,
  input  [31:0] io_fpu_store_data,
  input  [31:0] io_fpu_toint_data,
  output        io_fpu_dmem_resp_val,
  output [4:0]  io_fpu_dmem_resp_tag,
  output [31:0] io_fpu_dmem_resp_data,
  output        io_fpu_valid,
  input         io_fpu_fcsr_rdy,
  input         io_fpu_nack_mem,
  input         io_fpu_illegal_rm,
  output        io_fpu_killx,
  output        io_fpu_killm,
  input         io_fpu_dec_wen,
  input         io_fpu_dec_ren1,
  input         io_fpu_dec_ren2,
  input         io_fpu_dec_ren3,
  input         io_fpu_sboard_set,
  input         io_fpu_sboard_clr,
  input  [4:0]  io_fpu_sboard_clra,
  output        io_rocc_cmd_valid,
  output        io_wfi
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
`endif // RANDOMIZE_REG_INIT
  wire  ibuf_clock;
  wire  ibuf_reset;
  wire  ibuf_io_imem_ready;
  wire  ibuf_io_imem_valid;
  wire  ibuf_io_imem_bits_btb_taken;
  wire  ibuf_io_imem_bits_btb_bridx;
  wire [4:0] ibuf_io_imem_bits_btb_entry;
  wire [7:0] ibuf_io_imem_bits_btb_bht_history;
  wire [31:0] ibuf_io_imem_bits_pc;
  wire [31:0] ibuf_io_imem_bits_data;
  wire  ibuf_io_imem_bits_xcpt_pf_inst;
  wire  ibuf_io_imem_bits_xcpt_ae_inst;
  wire  ibuf_io_imem_bits_replay;
  wire  ibuf_io_kill;
  wire [31:0] ibuf_io_pc;
  wire [4:0] ibuf_io_btb_resp_entry;
  wire [7:0] ibuf_io_btb_resp_bht_history;
  wire  ibuf_io_inst_0_ready;
  wire  ibuf_io_inst_0_valid;
  wire  ibuf_io_inst_0_bits_xcpt0_pf_inst;
  wire  ibuf_io_inst_0_bits_xcpt0_ae_inst;
  wire  ibuf_io_inst_0_bits_xcpt1_pf_inst;
  wire  ibuf_io_inst_0_bits_xcpt1_gf_inst;
  wire  ibuf_io_inst_0_bits_xcpt1_ae_inst;
  wire  ibuf_io_inst_0_bits_replay;
  wire  ibuf_io_inst_0_bits_rvc;
  wire [31:0] ibuf_io_inst_0_bits_inst_bits;
  wire [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs3;
  wire [31:0] ibuf_io_inst_0_bits_raw;
  reg [31:0] rf [0:30];
  wire  rf_id_rs_MPORT_en;
  wire [4:0] rf_id_rs_MPORT_addr;
  wire [31:0] rf_id_rs_MPORT_data;
  wire  rf_id_rs_MPORT_1_en;
  wire [4:0] rf_id_rs_MPORT_1_addr;
  wire [31:0] rf_id_rs_MPORT_1_data;
  wire [31:0] rf_MPORT_data;
  wire [4:0] rf_MPORT_addr;
  wire  rf_MPORT_mask;
  wire  rf_MPORT_en;
  wire  csr_clock;
  wire  csr_reset;
  wire  csr_io_ungated_clock;
  wire  csr_io_interrupts_debug;
  wire  csr_io_interrupts_mtip;
  wire  csr_io_interrupts_msip;
  wire  csr_io_interrupts_meip;
  wire  csr_io_interrupts_seip;
  wire  csr_io_hartid;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [31:0] csr_io_rw_rdata;
  wire [31:0] csr_io_rw_wdata;
  wire [31:0] csr_io_decode_0_inst;
  wire  csr_io_decode_0_fp_illegal;
  wire  csr_io_decode_0_fp_csr;
  wire  csr_io_decode_0_rocc_illegal;
  wire  csr_io_decode_0_read_illegal;
  wire  csr_io_decode_0_write_illegal;
  wire  csr_io_decode_0_write_flush;
  wire  csr_io_decode_0_system_illegal;
  wire  csr_io_csr_stall;
  wire  csr_io_eret;
  wire  csr_io_singleStep;
  wire  csr_io_status_debug;
  wire  csr_io_status_cease;
  wire  csr_io_status_wfi;
  wire [31:0] csr_io_status_isa;
  wire [1:0] csr_io_status_dprv;
  wire  csr_io_status_dv;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_v;
  wire  csr_io_status_sd;
  wire [22:0] csr_io_status_zero2;
  wire  csr_io_status_mpv;
  wire  csr_io_status_gva;
  wire  csr_io_status_mbe;
  wire  csr_io_status_sbe;
  wire [1:0] csr_io_status_sxl;
  wire [1:0] csr_io_status_uxl;
  wire  csr_io_status_sd_rv32;
  wire [7:0] csr_io_status_zero1;
  wire  csr_io_status_tsr;
  wire  csr_io_status_tw;
  wire  csr_io_status_tvm;
  wire  csr_io_status_mxr;
  wire  csr_io_status_sum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_vs;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_ube;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire  csr_io_ptbr_mode;
  wire [21:0] csr_io_ptbr_ppn;
  wire [31:0] csr_io_evec;
  wire  csr_io_exception;
  wire  csr_io_retire;
  wire [31:0] csr_io_cause;
  wire [31:0] csr_io_pc;
  wire [31:0] csr_io_tval;
  wire  csr_io_gva;
  wire [31:0] csr_io_time;
  wire [2:0] csr_io_fcsr_rm;
  wire  csr_io_fcsr_flags_valid;
  wire [4:0] csr_io_fcsr_flags_bits;
  wire  csr_io_interrupt;
  wire [31:0] csr_io_interrupt_cause;
  wire  csr_io_bp_0_control_action;
  wire [1:0] csr_io_bp_0_control_tmatch;
  wire  csr_io_bp_0_control_m;
  wire  csr_io_bp_0_control_s;
  wire  csr_io_bp_0_control_u;
  wire  csr_io_bp_0_control_x;
  wire  csr_io_bp_0_control_w;
  wire  csr_io_bp_0_control_r;
  wire [31:0] csr_io_bp_0_address;
  wire  csr_io_pmp_0_cfg_l;
  wire [1:0] csr_io_pmp_0_cfg_a;
  wire  csr_io_pmp_0_cfg_x;
  wire  csr_io_pmp_0_cfg_w;
  wire  csr_io_pmp_0_cfg_r;
  wire [29:0] csr_io_pmp_0_addr;
  wire [31:0] csr_io_pmp_0_mask;
  wire  csr_io_pmp_1_cfg_l;
  wire [1:0] csr_io_pmp_1_cfg_a;
  wire  csr_io_pmp_1_cfg_x;
  wire  csr_io_pmp_1_cfg_w;
  wire  csr_io_pmp_1_cfg_r;
  wire [29:0] csr_io_pmp_1_addr;
  wire [31:0] csr_io_pmp_1_mask;
  wire  csr_io_pmp_2_cfg_l;
  wire [1:0] csr_io_pmp_2_cfg_a;
  wire  csr_io_pmp_2_cfg_x;
  wire  csr_io_pmp_2_cfg_w;
  wire  csr_io_pmp_2_cfg_r;
  wire [29:0] csr_io_pmp_2_addr;
  wire [31:0] csr_io_pmp_2_mask;
  wire  csr_io_pmp_3_cfg_l;
  wire [1:0] csr_io_pmp_3_cfg_a;
  wire  csr_io_pmp_3_cfg_x;
  wire  csr_io_pmp_3_cfg_w;
  wire  csr_io_pmp_3_cfg_r;
  wire [29:0] csr_io_pmp_3_addr;
  wire [31:0] csr_io_pmp_3_mask;
  wire  csr_io_pmp_4_cfg_l;
  wire [1:0] csr_io_pmp_4_cfg_a;
  wire  csr_io_pmp_4_cfg_x;
  wire  csr_io_pmp_4_cfg_w;
  wire  csr_io_pmp_4_cfg_r;
  wire [29:0] csr_io_pmp_4_addr;
  wire [31:0] csr_io_pmp_4_mask;
  wire  csr_io_pmp_5_cfg_l;
  wire [1:0] csr_io_pmp_5_cfg_a;
  wire  csr_io_pmp_5_cfg_x;
  wire  csr_io_pmp_5_cfg_w;
  wire  csr_io_pmp_5_cfg_r;
  wire [29:0] csr_io_pmp_5_addr;
  wire [31:0] csr_io_pmp_5_mask;
  wire  csr_io_pmp_6_cfg_l;
  wire [1:0] csr_io_pmp_6_cfg_a;
  wire  csr_io_pmp_6_cfg_x;
  wire  csr_io_pmp_6_cfg_w;
  wire  csr_io_pmp_6_cfg_r;
  wire [29:0] csr_io_pmp_6_addr;
  wire [31:0] csr_io_pmp_6_mask;
  wire  csr_io_pmp_7_cfg_l;
  wire [1:0] csr_io_pmp_7_cfg_a;
  wire  csr_io_pmp_7_cfg_x;
  wire  csr_io_pmp_7_cfg_w;
  wire  csr_io_pmp_7_cfg_r;
  wire [29:0] csr_io_pmp_7_addr;
  wire [31:0] csr_io_pmp_7_mask;
  wire  csr_io_inhibit_cycle;
  wire [31:0] csr_io_inst_0;
  wire  csr_io_trace_0_valid;
  wire [31:0] csr_io_trace_0_iaddr;
  wire [31:0] csr_io_trace_0_insn;
  wire  csr_io_trace_0_exception;
  wire [31:0] csr_io_customCSRs_0_value;
  wire  bpu_io_status_debug;
  wire [1:0] bpu_io_status_prv;
  wire  bpu_io_bp_0_control_action;
  wire [1:0] bpu_io_bp_0_control_tmatch;
  wire  bpu_io_bp_0_control_m;
  wire  bpu_io_bp_0_control_s;
  wire  bpu_io_bp_0_control_u;
  wire  bpu_io_bp_0_control_x;
  wire  bpu_io_bp_0_control_w;
  wire  bpu_io_bp_0_control_r;
  wire [31:0] bpu_io_bp_0_address;
  wire [31:0] bpu_io_pc;
  wire [31:0] bpu_io_ea;
  wire  bpu_io_xcpt_if;
  wire  bpu_io_xcpt_ld;
  wire  bpu_io_xcpt_st;
  wire  bpu_io_debug_if;
  wire  bpu_io_debug_ld;
  wire  bpu_io_debug_st;
  wire [3:0] alu_io_fn;
  wire [31:0] alu_io_in2;
  wire [31:0] alu_io_in1;
  wire [31:0] alu_io_out;
  wire [31:0] alu_io_adder_out;
  wire  alu_io_cmp_out;
  wire  div_clock;
  wire  div_reset;
  wire  div_io_req_ready;
  wire  div_io_req_valid;
  wire [3:0] div_io_req_bits_fn;
  wire [31:0] div_io_req_bits_in1;
  wire [31:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire  div_io_kill;
  wire  div_io_resp_ready;
  wire  div_io_resp_valid;
  wire [31:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire  PlusArgTimeout_clock;
  wire  PlusArgTimeout_reset;
  wire [31:0] PlusArgTimeout_io_count;
  reg  id_reg_pause;
  reg  imem_might_request_reg;
  reg  ex_ctrl_fp;
  reg  ex_ctrl_rocc;
  reg  ex_ctrl_branch;
  reg  ex_ctrl_jal;
  reg  ex_ctrl_jalr;
  reg  ex_ctrl_rxs2;
  reg  ex_ctrl_rxs1;
  reg [1:0] ex_ctrl_sel_alu2;
  reg [1:0] ex_ctrl_sel_alu1;
  reg [2:0] ex_ctrl_sel_imm;
  reg [3:0] ex_ctrl_alu_fn;
  reg  ex_ctrl_mem;
  reg [4:0] ex_ctrl_mem_cmd;
  reg  ex_ctrl_rfs1;
  reg  ex_ctrl_rfs2;
  reg  ex_ctrl_wfd;
  reg  ex_ctrl_mul;
  reg  ex_ctrl_div;
  reg  ex_ctrl_wxd;
  reg [2:0] ex_ctrl_csr;
  reg  ex_ctrl_fence_i;
  reg  mem_ctrl_fp;
  reg  mem_ctrl_rocc;
  reg  mem_ctrl_branch;
  reg  mem_ctrl_jal;
  reg  mem_ctrl_jalr;
  reg  mem_ctrl_rxs2;
  reg  mem_ctrl_rxs1;
  reg  mem_ctrl_mem;
  reg  mem_ctrl_rfs1;
  reg  mem_ctrl_rfs2;
  reg  mem_ctrl_wfd;
  reg  mem_ctrl_mul;
  reg  mem_ctrl_div;
  reg  mem_ctrl_wxd;
  reg [2:0] mem_ctrl_csr;
  reg  mem_ctrl_fence_i;
  reg  wb_ctrl_rocc;
  reg  wb_ctrl_rxs2;
  reg  wb_ctrl_rxs1;
  reg  wb_ctrl_mem;
  reg  wb_ctrl_rfs1;
  reg  wb_ctrl_rfs2;
  reg  wb_ctrl_wfd;
  reg  wb_ctrl_div;
  reg  wb_ctrl_wxd;
  reg [2:0] wb_ctrl_csr;
  reg  wb_ctrl_fence_i;
  reg  ex_reg_xcpt_interrupt;
  reg  ex_reg_valid;
  reg  ex_reg_rvc;
  reg [4:0] ex_reg_btb_resp_entry;
  reg [7:0] ex_reg_btb_resp_bht_history;
  reg  ex_reg_xcpt;
  reg  ex_reg_flush_pipe;
  reg  ex_reg_load_use;
  reg [31:0] ex_reg_cause;
  reg  ex_reg_replay;
  reg [31:0] ex_reg_pc;
  reg [1:0] ex_reg_mem_size;
  reg [31:0] ex_reg_inst;
  reg [31:0] ex_reg_raw_inst;
  reg  mem_reg_xcpt_interrupt;
  reg  mem_reg_valid;
  reg  mem_reg_rvc;
  reg [4:0] mem_reg_btb_resp_entry;
  reg [7:0] mem_reg_btb_resp_bht_history;
  reg  mem_reg_xcpt;
  reg  mem_reg_replay;
  reg  mem_reg_flush_pipe;
  reg [31:0] mem_reg_cause;
  reg  mem_reg_slow_bypass;
  reg  mem_reg_load;
  reg  mem_reg_store;
  reg  mem_reg_sfence;
  reg [31:0] mem_reg_pc;
  reg [31:0] mem_reg_inst;
  reg [1:0] mem_reg_mem_size;
  reg  mem_reg_hls_or_dv;
  reg [31:0] mem_reg_raw_inst;
  reg [31:0] mem_reg_wdata;
  reg [31:0] mem_reg_rs2;
  reg  mem_br_taken;
  reg  wb_reg_valid;
  reg  wb_reg_xcpt;
  reg  wb_reg_replay;
  reg  wb_reg_flush_pipe;
  reg [31:0] wb_reg_cause;
  reg  wb_reg_sfence;
  reg [31:0] wb_reg_pc;
  reg [1:0] wb_reg_mem_size;
  reg  wb_reg_hls_or_dv;
  reg [31:0] wb_reg_inst;
  reg [31:0] wb_reg_raw_inst;
  reg [31:0] wb_reg_wdata;
  wire  replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
  wire  replay_wb_rocc = wb_reg_valid & wb_ctrl_rocc;
  wire  replay_wb = replay_wb_common | replay_wb_rocc;
  wire  _T_96 = wb_reg_valid & wb_ctrl_mem;
  wire  _T_97 = wb_reg_valid & wb_ctrl_mem & io_dmem_s2_xcpt_pf_st;
  wire  _T_99 = _T_96 & io_dmem_s2_xcpt_pf_ld;
  wire  _T_105 = _T_96 & io_dmem_s2_xcpt_ae_st;
  wire  _T_107 = _T_96 & io_dmem_s2_xcpt_ae_ld;
  wire  _T_109 = _T_96 & io_dmem_s2_xcpt_ma_st;
  wire  _T_111 = _T_96 & io_dmem_s2_xcpt_ma_ld;
  wire  wb_xcpt = wb_reg_xcpt | _T_97 | _T_99 | _T_105 | _T_107 | _T_109 | _T_111;
  wire  take_pc_wb = replay_wb | wb_xcpt | csr_io_eret | wb_reg_flush_pipe;
  wire  _take_pc_mem_T = ~mem_reg_xcpt;
  wire  ex_pc_valid = ex_reg_valid | ex_reg_replay | ex_reg_xcpt_interrupt;
  wire  _mem_br_target_T_1 = mem_ctrl_branch & mem_br_taken;
  wire  mem_br_target_sign = mem_reg_inst[31];
  wire  mem_br_target_hi_hi_hi = mem_reg_inst[31];
  wire [10:0] mem_br_target_hi_hi_lo = {11{mem_br_target_sign}};
  wire [7:0] mem_br_target_hi_lo_hi = {8{mem_br_target_sign}};
  wire  mem_br_target_hi_lo_lo = mem_reg_inst[7];
  wire [5:0] mem_br_target_b10_5 = mem_reg_inst[30:25];
  wire [3:0] mem_br_target_b4_1 = mem_reg_inst[11:8];
  wire [31:0] _mem_br_target_T_3 = {mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi,
    mem_br_target_hi_lo_lo,mem_br_target_b10_5,mem_br_target_b4_1,1'h0};
  wire [7:0] mem_br_target_hi_lo_hi_1 = mem_reg_inst[19:12];
  wire  mem_br_target_hi_lo_lo_1 = mem_reg_inst[20];
  wire [31:0] _mem_br_target_T_5 = {mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi_1,
    mem_br_target_hi_lo_lo_1,mem_br_target_b10_5,mem_reg_inst[24:21],1'h0};
  wire [3:0] _mem_br_target_T_6 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  wire [31:0] _mem_br_target_T_7 = mem_ctrl_jal ? $signed(_mem_br_target_T_5) : $signed({{28{_mem_br_target_T_6[3]}},
    _mem_br_target_T_6});
  wire [31:0] _mem_br_target_T_8 = mem_ctrl_branch & mem_br_taken ? $signed(_mem_br_target_T_3) : $signed(
    _mem_br_target_T_7);
  wire [31:0] mem_br_target = $signed(mem_reg_pc) + $signed(_mem_br_target_T_8);
  wire [31:0] _mem_npc_T_2 = mem_ctrl_jalr | mem_reg_sfence ? $signed(mem_reg_wdata) : $signed(mem_br_target);
  wire [31:0] mem_npc = $signed(_mem_npc_T_2) & -32'sh2;
  wire  _mem_wrong_npc_T_3 = ibuf_io_inst_0_valid | ibuf_io_imem_valid ? mem_npc != ibuf_io_pc : 1'h1;
  wire  mem_wrong_npc = ex_pc_valid ? mem_npc != ex_reg_pc : _mem_wrong_npc_T_3;
  wire  take_pc_mem = mem_reg_valid & ~mem_reg_xcpt & (mem_wrong_npc | mem_reg_sfence);
  wire  take_pc_mem_wb = take_pc_wb | take_pc_mem;
  wire [31:0] id_ctrl_decoder_decoded_plaInput = ibuf_io_inst_0_bits_inst_bits;
  wire [31:0] id_ctrl_decoder_decoded_invInputs = ~id_ctrl_decoder_decoded_plaInput;
  wire  id_ctrl_decoder_decoded_andMatrixInput_0 = id_ctrl_decoder_decoded_plaInput[0];
  wire  id_ctrl_decoder_decoded_andMatrixInput_1 = id_ctrl_decoder_decoded_plaInput[1];
  wire  id_ctrl_decoder_decoded_andMatrixInput_2 = id_ctrl_decoder_decoded_invInputs[2];
  wire  id_ctrl_decoder_decoded_andMatrixInput_3 = id_ctrl_decoder_decoded_invInputs[3];
  wire  id_ctrl_decoder_decoded_andMatrixInput_4 = id_ctrl_decoder_decoded_invInputs[4];
  wire  id_ctrl_decoder_decoded_andMatrixInput_5 = id_ctrl_decoder_decoded_invInputs[5];
  wire  id_ctrl_decoder_decoded_andMatrixInput_6 = id_ctrl_decoder_decoded_invInputs[6];
  wire  id_ctrl_decoder_decoded_andMatrixInput_7 = id_ctrl_decoder_decoded_invInputs[13];
  wire [7:0] _id_ctrl_decoder_decoded_T = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7};
  wire  _id_ctrl_decoder_decoded_T_1 = &_id_ctrl_decoder_decoded_T;
  wire  id_ctrl_decoder_decoded_andMatrixInput_6_1 = id_ctrl_decoder_decoded_invInputs[12];
  wire [7:0] _id_ctrl_decoder_decoded_T_2 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_7};
  wire  _id_ctrl_decoder_decoded_T_3 = &_id_ctrl_decoder_decoded_T_2;
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_2 = id_ctrl_decoder_decoded_invInputs[14];
  wire [7:0] _id_ctrl_decoder_decoded_T_4 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_5 = &_id_ctrl_decoder_decoded_T_4;
  wire [7:0] _id_ctrl_decoder_decoded_T_6 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_7 = &_id_ctrl_decoder_decoded_T_6;
  wire  id_ctrl_decoder_decoded_andMatrixInput_2_4 = id_ctrl_decoder_decoded_plaInput[2];
  wire  id_ctrl_decoder_decoded_andMatrixInput_3_4 = id_ctrl_decoder_decoded_plaInput[3];
  wire [8:0] _id_ctrl_decoder_decoded_T_8 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_9 = &_id_ctrl_decoder_decoded_T_8;
  wire  id_ctrl_decoder_decoded_andMatrixInput_4_5 = id_ctrl_decoder_decoded_plaInput[4];
  wire [5:0] _id_ctrl_decoder_decoded_T_10 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_6};
  wire  _id_ctrl_decoder_decoded_T_11 = &_id_ctrl_decoder_decoded_T_10;
  wire [6:0] _id_ctrl_decoder_decoded_T_12 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6};
  wire  _id_ctrl_decoder_decoded_T_13 = &_id_ctrl_decoder_decoded_T_12;
  wire  id_ctrl_decoder_decoded_andMatrixInput_5_7 = id_ctrl_decoder_decoded_plaInput[5];
  wire [8:0] _id_ctrl_decoder_decoded_T_14 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_15 = &_id_ctrl_decoder_decoded_T_14;
  wire [7:0] _id_ctrl_decoder_decoded_T_16 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_17 = &_id_ctrl_decoder_decoded_T_16;
  wire [8:0] _id_ctrl_decoder_decoded_T_18 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_19 = &_id_ctrl_decoder_decoded_T_18;
  wire  id_ctrl_decoder_decoded_andMatrixInput_10 = id_ctrl_decoder_decoded_invInputs[25];
  wire  id_ctrl_decoder_decoded_andMatrixInput_11 = id_ctrl_decoder_decoded_invInputs[26];
  wire  id_ctrl_decoder_decoded_andMatrixInput_12 = id_ctrl_decoder_decoded_invInputs[27];
  wire  id_ctrl_decoder_decoded_andMatrixInput_13 = id_ctrl_decoder_decoded_invInputs[28];
  wire  id_ctrl_decoder_decoded_andMatrixInput_14 = id_ctrl_decoder_decoded_invInputs[29];
  wire  id_ctrl_decoder_decoded_andMatrixInput_15 = id_ctrl_decoder_decoded_invInputs[31];
  wire [7:0] id_ctrl_decoder_decoded_lo_10 = {id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] _id_ctrl_decoder_decoded_T_20 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_lo_10};
  wire  _id_ctrl_decoder_decoded_T_21 = &_id_ctrl_decoder_decoded_T_20;
  wire  id_ctrl_decoder_decoded_andMatrixInput_11_1 = id_ctrl_decoder_decoded_invInputs[30];
  wire [5:0] id_ctrl_decoder_decoded_lo_11 = {id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [12:0] _id_ctrl_decoder_decoded_T_22 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_11};
  wire  _id_ctrl_decoder_decoded_T_23 = &_id_ctrl_decoder_decoded_T_22;
  wire  id_ctrl_decoder_decoded_andMatrixInput_4_12 = id_ctrl_decoder_decoded_plaInput[6];
  wire [4:0] _id_ctrl_decoder_decoded_T_24 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12};
  wire  _id_ctrl_decoder_decoded_T_25 = &_id_ctrl_decoder_decoded_T_24;
  wire [6:0] _id_ctrl_decoder_decoded_T_26 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11};
  wire  _id_ctrl_decoder_decoded_T_27 = &_id_ctrl_decoder_decoded_T_26;
  wire [5:0] id_ctrl_decoder_decoded_lo_14 = {id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [11:0] _id_ctrl_decoder_decoded_T_28 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_lo_14};
  wire  _id_ctrl_decoder_decoded_T_29 = &_id_ctrl_decoder_decoded_T_28;
  wire [7:0] _id_ctrl_decoder_decoded_T_30 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7};
  wire  _id_ctrl_decoder_decoded_T_31 = &_id_ctrl_decoder_decoded_T_30;
  wire [8:0] _id_ctrl_decoder_decoded_T_32 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_33 = &_id_ctrl_decoder_decoded_T_32;
  wire [8:0] _id_ctrl_decoder_decoded_T_34 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_3,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_35 = &_id_ctrl_decoder_decoded_T_34;
  wire [9:0] _id_ctrl_decoder_decoded_T_36 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_37 = &_id_ctrl_decoder_decoded_T_36;
  wire [6:0] _id_ctrl_decoder_decoded_T_38 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12};
  wire  _id_ctrl_decoder_decoded_T_39 = &_id_ctrl_decoder_decoded_T_38;
  wire  id_ctrl_decoder_decoded_andMatrixInput_4_20 = id_ctrl_decoder_decoded_invInputs[7];
  wire  id_ctrl_decoder_decoded_andMatrixInput_5_19 = id_ctrl_decoder_decoded_invInputs[8];
  wire  id_ctrl_decoder_decoded_andMatrixInput_6_18 = id_ctrl_decoder_decoded_invInputs[9];
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_15 = id_ctrl_decoder_decoded_invInputs[10];
  wire  id_ctrl_decoder_decoded_andMatrixInput_8_9 = id_ctrl_decoder_decoded_invInputs[11];
  wire  id_ctrl_decoder_decoded_andMatrixInput_12_2 = id_ctrl_decoder_decoded_invInputs[15];
  wire  id_ctrl_decoder_decoded_andMatrixInput_13_1 = id_ctrl_decoder_decoded_invInputs[16];
  wire  id_ctrl_decoder_decoded_andMatrixInput_14_1 = id_ctrl_decoder_decoded_invInputs[17];
  wire  id_ctrl_decoder_decoded_andMatrixInput_15_1 = id_ctrl_decoder_decoded_invInputs[18];
  wire  id_ctrl_decoder_decoded_andMatrixInput_16 = id_ctrl_decoder_decoded_invInputs[19];
  wire  id_ctrl_decoder_decoded_andMatrixInput_17 = id_ctrl_decoder_decoded_invInputs[21];
  wire  id_ctrl_decoder_decoded_andMatrixInput_18 = id_ctrl_decoder_decoded_invInputs[22];
  wire  id_ctrl_decoder_decoded_andMatrixInput_19 = id_ctrl_decoder_decoded_invInputs[23];
  wire  id_ctrl_decoder_decoded_andMatrixInput_20 = id_ctrl_decoder_decoded_invInputs[24];
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_15 = {id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [13:0] id_ctrl_decoder_decoded_lo_20 = {id_ctrl_decoder_decoded_andMatrixInput_14_1,
    id_ctrl_decoder_decoded_andMatrixInput_15_1,id_ctrl_decoder_decoded_andMatrixInput_16,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_lo_lo_15
    };
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_18 = {id_ctrl_decoder_decoded_andMatrixInput_7_15,
    id_ctrl_decoder_decoded_andMatrixInput_8_9,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_12_2,id_ctrl_decoder_decoded_andMatrixInput_13_1};
  wire [27:0] _id_ctrl_decoder_decoded_T_40 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_4_5,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_4_20,
    id_ctrl_decoder_decoded_andMatrixInput_5_19,id_ctrl_decoder_decoded_andMatrixInput_6_18,
    id_ctrl_decoder_decoded_hi_lo_18,id_ctrl_decoder_decoded_lo_20};
  wire  _id_ctrl_decoder_decoded_T_41 = &_id_ctrl_decoder_decoded_T_40;
  wire [14:0] id_ctrl_decoder_decoded_lo_21 = {id_ctrl_decoder_decoded_andMatrixInput_13_1,
    id_ctrl_decoder_decoded_andMatrixInput_14_1,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_17,
    id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_lo_lo_15};
  wire [7:0] id_ctrl_decoder_decoded_hi_lo_19 = {id_ctrl_decoder_decoded_andMatrixInput_5_19,
    id_ctrl_decoder_decoded_andMatrixInput_6_18,id_ctrl_decoder_decoded_andMatrixInput_7_15,
    id_ctrl_decoder_decoded_andMatrixInput_8_9,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_12_2};
  wire [30:0] _id_ctrl_decoder_decoded_T_42 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_hi_lo_19,id_ctrl_decoder_decoded_lo_21};
  wire  _id_ctrl_decoder_decoded_T_43 = &_id_ctrl_decoder_decoded_T_42;
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_17 = id_ctrl_decoder_decoded_plaInput[12];
  wire [9:0] _id_ctrl_decoder_decoded_T_44 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_45 = &_id_ctrl_decoder_decoded_T_44;
  wire [14:0] _id_ctrl_decoder_decoded_T_46 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_lo_15};
  wire  _id_ctrl_decoder_decoded_T_47 = &_id_ctrl_decoder_decoded_T_46;
  wire [7:0] id_ctrl_decoder_decoded_lo_24 = {id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] _id_ctrl_decoder_decoded_T_48 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_lo_24};
  wire  _id_ctrl_decoder_decoded_T_49 = &_id_ctrl_decoder_decoded_T_48;
  wire [7:0] _id_ctrl_decoder_decoded_T_50 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_7};
  wire  _id_ctrl_decoder_decoded_T_51 = &_id_ctrl_decoder_decoded_T_50;
  wire [8:0] _id_ctrl_decoder_decoded_T_52 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_andMatrixInput_7};
  wire  _id_ctrl_decoder_decoded_T_53 = &_id_ctrl_decoder_decoded_T_52;
  wire [8:0] _id_ctrl_decoder_decoded_T_54 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_55 = &_id_ctrl_decoder_decoded_T_54;
  wire [7:0] _id_ctrl_decoder_decoded_T_56 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7_17};
  wire  _id_ctrl_decoder_decoded_T_57 = &_id_ctrl_decoder_decoded_T_56;
  wire  id_ctrl_decoder_decoded_andMatrixInput_6_27 = id_ctrl_decoder_decoded_plaInput[13];
  wire [7:0] _id_ctrl_decoder_decoded_T_58 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_3,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_59 = &_id_ctrl_decoder_decoded_T_58;
  wire [8:0] _id_ctrl_decoder_decoded_T_60 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_3,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_61 = &_id_ctrl_decoder_decoded_T_60;
  wire [8:0] _id_ctrl_decoder_decoded_T_62 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_63 = &_id_ctrl_decoder_decoded_T_62;
  wire [9:0] _id_ctrl_decoder_decoded_T_64 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_65 = &_id_ctrl_decoder_decoded_T_64;
  wire [7:0] _id_ctrl_decoder_decoded_T_66 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_27};
  wire  _id_ctrl_decoder_decoded_T_67 = &_id_ctrl_decoder_decoded_T_66;
  wire [8:0] _id_ctrl_decoder_decoded_T_68 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_69 = &_id_ctrl_decoder_decoded_T_68;
  wire [8:0] _id_ctrl_decoder_decoded_T_70 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_3,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_71 = &_id_ctrl_decoder_decoded_T_70;
  wire [9:0] _id_ctrl_decoder_decoded_T_72 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_73 = &_id_ctrl_decoder_decoded_T_72;
  wire [5:0] id_ctrl_decoder_decoded_lo_37 = {id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_7_2,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13};
  wire [11:0] _id_ctrl_decoder_decoded_T_74 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_lo_37};
  wire  _id_ctrl_decoder_decoded_T_75 = &_id_ctrl_decoder_decoded_T_74;
  wire [14:0] _id_ctrl_decoder_decoded_T_76 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_lo_lo_15};
  wire  _id_ctrl_decoder_decoded_T_77 = &_id_ctrl_decoder_decoded_T_76;
  wire [7:0] id_ctrl_decoder_decoded_lo_39 = {id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] _id_ctrl_decoder_decoded_T_78 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_lo_39};
  wire  _id_ctrl_decoder_decoded_T_79 = &_id_ctrl_decoder_decoded_T_78;
  wire [7:0] _id_ctrl_decoder_decoded_T_80 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_27};
  wire  _id_ctrl_decoder_decoded_T_81 = &_id_ctrl_decoder_decoded_T_80;
  wire [8:0] _id_ctrl_decoder_decoded_T_82 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire  _id_ctrl_decoder_decoded_T_83 = &_id_ctrl_decoder_decoded_T_82;
  wire [8:0] _id_ctrl_decoder_decoded_T_84 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_andMatrixInput_6_27};
  wire  _id_ctrl_decoder_decoded_T_85 = &_id_ctrl_decoder_decoded_T_84;
  wire [6:0] id_ctrl_decoder_decoded_lo_43 = {id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [14:0] _id_ctrl_decoder_decoded_T_86 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_lo_43};
  wire  _id_ctrl_decoder_decoded_T_87 = &_id_ctrl_decoder_decoded_T_86;
  wire  id_ctrl_decoder_decoded_andMatrixInput_8_28 = id_ctrl_decoder_decoded_plaInput[14];
  wire [8:0] _id_ctrl_decoder_decoded_T_88 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_89 = &_id_ctrl_decoder_decoded_T_88;
  wire [6:0] id_ctrl_decoder_decoded_lo_45 = {id_ctrl_decoder_decoded_andMatrixInput_8_28,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [13:0] _id_ctrl_decoder_decoded_T_90 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_45};
  wire  _id_ctrl_decoder_decoded_T_91 = &_id_ctrl_decoder_decoded_T_90;
  wire [7:0] _id_ctrl_decoder_decoded_T_92 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_93 = &_id_ctrl_decoder_decoded_T_92;
  wire [6:0] id_ctrl_decoder_decoded_lo_47 = {id_ctrl_decoder_decoded_andMatrixInput_8_28,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [14:0] _id_ctrl_decoder_decoded_T_94 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_47};
  wire  _id_ctrl_decoder_decoded_T_95 = &_id_ctrl_decoder_decoded_T_94;
  wire [7:0] id_ctrl_decoder_decoded_lo_48 = {id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_8_28,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] _id_ctrl_decoder_decoded_T_96 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_lo_48};
  wire  _id_ctrl_decoder_decoded_T_97 = &_id_ctrl_decoder_decoded_T_96;
  wire [7:0] id_ctrl_decoder_decoded_lo_49 = {id_ctrl_decoder_decoded_andMatrixInput_8_28,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] _id_ctrl_decoder_decoded_T_98 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_49};
  wire  _id_ctrl_decoder_decoded_T_99 = &_id_ctrl_decoder_decoded_T_98;
  wire [15:0] _id_ctrl_decoder_decoded_T_100 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_lo_48};
  wire  _id_ctrl_decoder_decoded_T_101 = &_id_ctrl_decoder_decoded_T_100;
  wire [14:0] _id_ctrl_decoder_decoded_T_102 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_lo_45};
  wire  _id_ctrl_decoder_decoded_T_103 = &_id_ctrl_decoder_decoded_T_102;
  wire [7:0] _id_ctrl_decoder_decoded_T_104 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_105 = &_id_ctrl_decoder_decoded_T_104;
  wire [8:0] _id_ctrl_decoder_decoded_T_106 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_107 = &_id_ctrl_decoder_decoded_T_106;
  wire [8:0] _id_ctrl_decoder_decoded_T_108 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_109 = &_id_ctrl_decoder_decoded_T_108;
  wire [8:0] _id_ctrl_decoder_decoded_T_110 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_111 = &_id_ctrl_decoder_decoded_T_110;
  wire [14:0] _id_ctrl_decoder_decoded_T_112 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_lo_45};
  wire  _id_ctrl_decoder_decoded_T_113 = &_id_ctrl_decoder_decoded_T_112;
  wire [7:0] _id_ctrl_decoder_decoded_T_114 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_115 = &_id_ctrl_decoder_decoded_T_114;
  wire [8:0] _id_ctrl_decoder_decoded_T_116 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_117 = &_id_ctrl_decoder_decoded_T_116;
  wire [8:0] _id_ctrl_decoder_decoded_T_118 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_119 = &_id_ctrl_decoder_decoded_T_118;
  wire [9:0] _id_ctrl_decoder_decoded_T_120 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_8_28};
  wire  _id_ctrl_decoder_decoded_T_121 = &_id_ctrl_decoder_decoded_T_120;
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_56 = id_ctrl_decoder_decoded_plaInput[25];
  wire [6:0] id_ctrl_decoder_decoded_lo_61 = {id_ctrl_decoder_decoded_andMatrixInput_7_56,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [13:0] _id_ctrl_decoder_decoded_T_122 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_61};
  wire  _id_ctrl_decoder_decoded_T_123 = &_id_ctrl_decoder_decoded_T_122;
  wire [14:0] _id_ctrl_decoder_decoded_T_124 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_17,id_ctrl_decoder_decoded_lo_61};
  wire  _id_ctrl_decoder_decoded_T_125 = &_id_ctrl_decoder_decoded_T_124;
  wire [14:0] _id_ctrl_decoder_decoded_T_126 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_lo_61};
  wire  _id_ctrl_decoder_decoded_T_127 = &_id_ctrl_decoder_decoded_T_126;
  wire  id_ctrl_decoder_decoded_andMatrixInput_10_21 = id_ctrl_decoder_decoded_plaInput[27];
  wire [6:0] id_ctrl_decoder_decoded_lo_64 = {id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_10_21,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [13:0] _id_ctrl_decoder_decoded_T_128 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_64};
  wire  _id_ctrl_decoder_decoded_T_129 = &_id_ctrl_decoder_decoded_T_128;
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_60 = id_ctrl_decoder_decoded_invInputs[20];
  wire  id_ctrl_decoder_decoded_andMatrixInput_13_19 = id_ctrl_decoder_decoded_plaInput[28];
  wire [7:0] id_ctrl_decoder_decoded_lo_65 = {id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13_19,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [16:0] _id_ctrl_decoder_decoded_T_130 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_60,id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_lo_65}
    ;
  wire  _id_ctrl_decoder_decoded_T_131 = &_id_ctrl_decoder_decoded_T_130;
  wire [4:0] id_ctrl_decoder_decoded_lo_lo_61 = {id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13_19,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [9:0] id_ctrl_decoder_decoded_lo_66 = {id_ctrl_decoder_decoded_andMatrixInput_7_60,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13_19,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [9:0] id_ctrl_decoder_decoded_hi_66 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_7_2};
  wire [19:0] _id_ctrl_decoder_decoded_T_132 = {id_ctrl_decoder_decoded_hi_66,id_ctrl_decoder_decoded_lo_66};
  wire  _id_ctrl_decoder_decoded_T_133 = &_id_ctrl_decoder_decoded_T_132;
  wire  id_ctrl_decoder_decoded_andMatrixInput_18_3 = id_ctrl_decoder_decoded_plaInput[21];
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_62 = {id_ctrl_decoder_decoded_andMatrixInput_20,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13_19,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [13:0] id_ctrl_decoder_decoded_lo_67 = {id_ctrl_decoder_decoded_andMatrixInput_14_1,
    id_ctrl_decoder_decoded_andMatrixInput_15_1,id_ctrl_decoder_decoded_andMatrixInput_16,
    id_ctrl_decoder_decoded_andMatrixInput_7_60,id_ctrl_decoder_decoded_andMatrixInput_18_3,
    id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_62
    };
  wire [27:0] _id_ctrl_decoder_decoded_T_134 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_4_5,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_4_20,
    id_ctrl_decoder_decoded_andMatrixInput_5_19,id_ctrl_decoder_decoded_andMatrixInput_6_18,
    id_ctrl_decoder_decoded_hi_lo_18,id_ctrl_decoder_decoded_lo_67};
  wire  _id_ctrl_decoder_decoded_T_135 = &_id_ctrl_decoder_decoded_T_134;
  wire [14:0] id_ctrl_decoder_decoded_lo_68 = {id_ctrl_decoder_decoded_andMatrixInput_13_1,
    id_ctrl_decoder_decoded_andMatrixInput_14_1,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_7_60,
    id_ctrl_decoder_decoded_andMatrixInput_18_3,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_62};
  wire [30:0] _id_ctrl_decoder_decoded_T_136 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_hi_lo_19,id_ctrl_decoder_decoded_lo_68};
  wire  _id_ctrl_decoder_decoded_T_137 = &_id_ctrl_decoder_decoded_T_136;
  wire  id_ctrl_decoder_decoded_andMatrixInput_17_5 = id_ctrl_decoder_decoded_plaInput[20];
  wire  id_ctrl_decoder_decoded_andMatrixInput_19_5 = id_ctrl_decoder_decoded_plaInput[22];
  wire [13:0] id_ctrl_decoder_decoded_lo_69 = {id_ctrl_decoder_decoded_andMatrixInput_14_1,
    id_ctrl_decoder_decoded_andMatrixInput_15_1,id_ctrl_decoder_decoded_andMatrixInput_16,
    id_ctrl_decoder_decoded_andMatrixInput_17_5,id_ctrl_decoder_decoded_andMatrixInput_17,
    id_ctrl_decoder_decoded_andMatrixInput_19_5,id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_lo_lo_62};
  wire [27:0] _id_ctrl_decoder_decoded_T_138 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_4_5,id_ctrl_decoder_decoded_andMatrixInput_5_7,
    id_ctrl_decoder_decoded_andMatrixInput_4_12,id_ctrl_decoder_decoded_andMatrixInput_4_20,
    id_ctrl_decoder_decoded_andMatrixInput_5_19,id_ctrl_decoder_decoded_andMatrixInput_6_18,
    id_ctrl_decoder_decoded_hi_lo_18,id_ctrl_decoder_decoded_lo_69};
  wire  _id_ctrl_decoder_decoded_T_139 = &_id_ctrl_decoder_decoded_T_138;
  wire [14:0] id_ctrl_decoder_decoded_lo_70 = {id_ctrl_decoder_decoded_andMatrixInput_13_1,
    id_ctrl_decoder_decoded_andMatrixInput_14_1,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_17_5,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_19_5,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_62};
  wire [30:0] _id_ctrl_decoder_decoded_T_140 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_hi_lo_19,id_ctrl_decoder_decoded_lo_70};
  wire  _id_ctrl_decoder_decoded_T_141 = &_id_ctrl_decoder_decoded_T_140;
  wire [7:0] id_ctrl_decoder_decoded_lo_71 = {id_ctrl_decoder_decoded_andMatrixInput_6_18,
    id_ctrl_decoder_decoded_andMatrixInput_7_56,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13_19,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [16:0] _id_ctrl_decoder_decoded_T_142 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_andMatrixInput_5_19,
    id_ctrl_decoder_decoded_lo_71};
  wire  _id_ctrl_decoder_decoded_T_143 = &_id_ctrl_decoder_decoded_T_142;
  wire [8:0] id_ctrl_decoder_decoded_lo_72 = {id_ctrl_decoder_decoded_andMatrixInput_6_18,
    id_ctrl_decoder_decoded_andMatrixInput_7_2,id_ctrl_decoder_decoded_andMatrixInput_7_56,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13_19,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [17:0] _id_ctrl_decoder_decoded_T_144 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_andMatrixInput_5_19,
    id_ctrl_decoder_decoded_lo_72};
  wire  _id_ctrl_decoder_decoded_T_145 = &_id_ctrl_decoder_decoded_T_144;
  wire [9:0] id_ctrl_decoder_decoded_lo_73 = {id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_7_56,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13_19,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [9:0] id_ctrl_decoder_decoded_hi_73 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_andMatrixInput_5_19,
    id_ctrl_decoder_decoded_andMatrixInput_6_18};
  wire [19:0] _id_ctrl_decoder_decoded_T_146 = {id_ctrl_decoder_decoded_hi_73,id_ctrl_decoder_decoded_lo_73};
  wire  _id_ctrl_decoder_decoded_T_147 = &_id_ctrl_decoder_decoded_T_146;
  wire [10:0] id_ctrl_decoder_decoded_lo_74 = {id_ctrl_decoder_decoded_andMatrixInput_8_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2,id_ctrl_decoder_decoded_andMatrixInput_7_56,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_lo_lo_61};
  wire [4:0] id_ctrl_decoder_decoded_hi_lo_72 = {id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_andMatrixInput_5_19,
    id_ctrl_decoder_decoded_andMatrixInput_6_18,id_ctrl_decoder_decoded_andMatrixInput_7_15};
  wire [21:0] _id_ctrl_decoder_decoded_T_148 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_hi_lo_72,id_ctrl_decoder_decoded_lo_74};
  wire  _id_ctrl_decoder_decoded_T_149 = &_id_ctrl_decoder_decoded_T_148;
  wire [6:0] id_ctrl_decoder_decoded_lo_75 = {id_ctrl_decoder_decoded_andMatrixInput_6_27,
    id_ctrl_decoder_decoded_andMatrixInput_7_2,id_ctrl_decoder_decoded_andMatrixInput_10_21,
    id_ctrl_decoder_decoded_andMatrixInput_13_19,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [14:0] _id_ctrl_decoder_decoded_T_150 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_lo_75};
  wire  _id_ctrl_decoder_decoded_T_151 = &_id_ctrl_decoder_decoded_T_150;
  wire  id_ctrl_decoder_decoded_andMatrixInput_13_30 = id_ctrl_decoder_decoded_plaInput[29];
  wire [6:0] id_ctrl_decoder_decoded_lo_76 = {id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_11_1};
  wire [14:0] _id_ctrl_decoder_decoded_T_152 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_lo_76};
  wire  _id_ctrl_decoder_decoded_T_153 = &_id_ctrl_decoder_decoded_T_152;
  wire [14:0] _id_ctrl_decoder_decoded_T_154 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_76};
  wire  _id_ctrl_decoder_decoded_T_155 = &_id_ctrl_decoder_decoded_T_154;
  wire [6:0] id_ctrl_decoder_decoded_lo_78 = {id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_11_1,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [14:0] _id_ctrl_decoder_decoded_T_156 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_78};
  wire  _id_ctrl_decoder_decoded_T_157 = &_id_ctrl_decoder_decoded_T_156;
  wire [7:0] id_ctrl_decoder_decoded_lo_79 = {id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] _id_ctrl_decoder_decoded_T_158 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_lo_79};
  wire  _id_ctrl_decoder_decoded_T_159 = &_id_ctrl_decoder_decoded_T_158;
  wire [5:0] id_ctrl_decoder_decoded_lo_80 = {id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_13_30};
  wire [12:0] _id_ctrl_decoder_decoded_T_160 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_80};
  wire  _id_ctrl_decoder_decoded_T_161 = &_id_ctrl_decoder_decoded_T_160;
  wire  id_ctrl_decoder_decoded_andMatrixInput_15_19 = id_ctrl_decoder_decoded_plaInput[30];
  wire [7:0] id_ctrl_decoder_decoded_lo_81 = {id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_15_19,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [16:0] _id_ctrl_decoder_decoded_T_162 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_81};
  wire  _id_ctrl_decoder_decoded_T_163 = &_id_ctrl_decoder_decoded_T_162;
  wire [5:0] id_ctrl_decoder_decoded_lo_82 = {id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_15_19};
  wire [12:0] _id_ctrl_decoder_decoded_T_164 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_82};
  wire  _id_ctrl_decoder_decoded_T_165 = &_id_ctrl_decoder_decoded_T_164;
  wire [7:0] id_ctrl_decoder_decoded_lo_83 = {id_ctrl_decoder_decoded_andMatrixInput_8_28,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_15_19,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] _id_ctrl_decoder_decoded_T_166 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_83};
  wire  _id_ctrl_decoder_decoded_T_167 = &_id_ctrl_decoder_decoded_T_166;
  wire [9:0] id_ctrl_decoder_decoded_hi_84 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7_60,id_ctrl_decoder_decoded_andMatrixInput_17,
    id_ctrl_decoder_decoded_andMatrixInput_18};
  wire [18:0] _id_ctrl_decoder_decoded_T_168 = {id_ctrl_decoder_decoded_hi_84,id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_10_21,
    id_ctrl_decoder_decoded_andMatrixInput_13_19,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_15_19,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire  _id_ctrl_decoder_decoded_T_169 = &_id_ctrl_decoder_decoded_T_168;
  wire  id_ctrl_decoder_decoded_andMatrixInput_20_7 = id_ctrl_decoder_decoded_plaInput[24];
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_80 = {id_ctrl_decoder_decoded_andMatrixInput_7_56,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_10_21,
    id_ctrl_decoder_decoded_andMatrixInput_13_19,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_15_19,id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [13:0] id_ctrl_decoder_decoded_lo_85 = {id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_7_60,
    id_ctrl_decoder_decoded_andMatrixInput_18_3,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20_7,
    id_ctrl_decoder_decoded_lo_lo_80};
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_83 = {id_ctrl_decoder_decoded_andMatrixInput_8_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2,id_ctrl_decoder_decoded_andMatrixInput_12_2,
    id_ctrl_decoder_decoded_andMatrixInput_13_1,id_ctrl_decoder_decoded_andMatrixInput_14_1};
  wire [27:0] _id_ctrl_decoder_decoded_T_170 = {id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_andMatrixInput_5_19,
    id_ctrl_decoder_decoded_andMatrixInput_6_18,id_ctrl_decoder_decoded_andMatrixInput_7_15,
    id_ctrl_decoder_decoded_hi_lo_83,id_ctrl_decoder_decoded_lo_85};
  wire  _id_ctrl_decoder_decoded_T_171 = &_id_ctrl_decoder_decoded_T_170;
  wire [7:0] id_ctrl_decoder_decoded_lo_lo_81 = {id_ctrl_decoder_decoded_andMatrixInput_20_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_56,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_10_21,id_ctrl_decoder_decoded_andMatrixInput_13_19,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_15_19,
    id_ctrl_decoder_decoded_andMatrixInput_15};
  wire [15:0] id_ctrl_decoder_decoded_lo_86 = {id_ctrl_decoder_decoded_andMatrixInput_13_1,
    id_ctrl_decoder_decoded_andMatrixInput_14_1,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_7_60,
    id_ctrl_decoder_decoded_andMatrixInput_18_3,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_81};
  wire [31:0] _id_ctrl_decoder_decoded_T_172 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_4_20,id_ctrl_decoder_decoded_hi_lo_19,id_ctrl_decoder_decoded_lo_86};
  wire  _id_ctrl_decoder_decoded_T_173 = &_id_ctrl_decoder_decoded_T_172;
  wire  id_ctrl_decoder_decoded_andMatrixInput_12_42 = id_ctrl_decoder_decoded_plaInput[31];
  wire [5:0] id_ctrl_decoder_decoded_lo_87 = {id_ctrl_decoder_decoded_andMatrixInput_6_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_27,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [12:0] _id_ctrl_decoder_decoded_T_174 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_4,
    id_ctrl_decoder_decoded_andMatrixInput_3_4,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5_7,id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_87};
  wire  _id_ctrl_decoder_decoded_T_175 = &_id_ctrl_decoder_decoded_T_174;
  wire [7:0] id_ctrl_decoder_decoded_lo_88 = {id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_11_1,
    id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [15:0] _id_ctrl_decoder_decoded_T_176 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_lo_88};
  wire  _id_ctrl_decoder_decoded_T_177 = &_id_ctrl_decoder_decoded_T_176;
  wire [15:0] _id_ctrl_decoder_decoded_T_178 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_lo_88};
  wire  _id_ctrl_decoder_decoded_T_179 = &_id_ctrl_decoder_decoded_T_178;
  wire [7:0] id_ctrl_decoder_decoded_lo_90 = {id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_14,id_ctrl_decoder_decoded_andMatrixInput_15_19,
    id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [16:0] _id_ctrl_decoder_decoded_T_180 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_lo_90};
  wire  _id_ctrl_decoder_decoded_T_181 = &_id_ctrl_decoder_decoded_T_180;
  wire [8:0] id_ctrl_decoder_decoded_lo_91 = {id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_15_19,id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [17:0] _id_ctrl_decoder_decoded_T_182 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_lo_91};
  wire  _id_ctrl_decoder_decoded_T_183 = &_id_ctrl_decoder_decoded_T_182;
  wire [8:0] id_ctrl_decoder_decoded_lo_92 = {id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13_19,id_ctrl_decoder_decoded_andMatrixInput_14,
    id_ctrl_decoder_decoded_andMatrixInput_15_19,id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [17:0] _id_ctrl_decoder_decoded_T_184 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_lo_92};
  wire  _id_ctrl_decoder_decoded_T_185 = &_id_ctrl_decoder_decoded_T_184;
  wire [9:0] id_ctrl_decoder_decoded_lo_93 = {id_ctrl_decoder_decoded_andMatrixInput_17,
    id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_15_19,
    id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [4:0] id_ctrl_decoder_decoded_hi_lo_91 = {id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_6_1,id_ctrl_decoder_decoded_andMatrixInput_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_2,id_ctrl_decoder_decoded_andMatrixInput_7_60};
  wire [20:0] _id_ctrl_decoder_decoded_T_186 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_hi_lo_91,id_ctrl_decoder_decoded_lo_93};
  wire  _id_ctrl_decoder_decoded_T_187 = &_id_ctrl_decoder_decoded_T_186;
  wire [9:0] id_ctrl_decoder_decoded_lo_94 = {id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_15_19,
    id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [4:0] id_ctrl_decoder_decoded_hi_lo_92 = {id_ctrl_decoder_decoded_andMatrixInput_4_12,
    id_ctrl_decoder_decoded_andMatrixInput_7,id_ctrl_decoder_decoded_andMatrixInput_7_2,
    id_ctrl_decoder_decoded_andMatrixInput_7_60,id_ctrl_decoder_decoded_andMatrixInput_17};
  wire [20:0] _id_ctrl_decoder_decoded_T_188 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_hi_lo_92,id_ctrl_decoder_decoded_lo_94};
  wire  _id_ctrl_decoder_decoded_T_189 = &_id_ctrl_decoder_decoded_T_188;
  wire [4:0] id_ctrl_decoder_decoded_lo_lo_90 = {id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13_19,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_15_19,id_ctrl_decoder_decoded_andMatrixInput_12_42};
  wire [10:0] id_ctrl_decoder_decoded_lo_95 = {id_ctrl_decoder_decoded_andMatrixInput_17,
    id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_lo_lo_90};
  wire [21:0] _id_ctrl_decoder_decoded_T_190 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_5,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_hi_lo_91,id_ctrl_decoder_decoded_lo_95};
  wire  _id_ctrl_decoder_decoded_T_191 = &_id_ctrl_decoder_decoded_T_190;
  wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T = {_id_ctrl_decoder_decoded_T_75,_id_ctrl_decoder_decoded_T_129,
    _id_ctrl_decoder_decoded_T_131};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_1 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_2 = |_id_ctrl_decoder_decoded_T_9;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_3 = |_id_ctrl_decoder_decoded_T_45;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_4 = |_id_ctrl_decoder_decoded_T_57;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_5 = |_id_ctrl_decoder_decoded_T_81;
  wire [6:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_6 = {_id_ctrl_decoder_decoded_T_41,_id_ctrl_decoder_decoded_T_57
    ,_id_ctrl_decoder_decoded_T_81,_id_ctrl_decoder_decoded_T_135,_id_ctrl_decoder_decoded_T_139,
    _id_ctrl_decoder_decoded_T_143,_id_ctrl_decoder_decoded_T_171};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_7 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_6;
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_1 = {_id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_75
    ,_id_ctrl_decoder_decoded_T_81,_id_ctrl_decoder_decoded_T_95,_id_ctrl_decoder_decoded_T_129,
    _id_ctrl_decoder_decoded_T_131,_id_ctrl_decoder_decoded_T_177,_id_ctrl_decoder_decoded_T_179,
    _id_ctrl_decoder_decoded_T_183,_id_ctrl_decoder_decoded_T_189};
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_2 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_3,
    _id_ctrl_decoder_decoded_T_5,_id_ctrl_decoder_decoded_T_11,_id_ctrl_decoder_decoded_T_21,
    _id_ctrl_decoder_decoded_T_23,_id_ctrl_decoder_decoded_T_37,_id_ctrl_decoder_decoded_T_39,
    _id_ctrl_decoder_decoded_T_47,_id_ctrl_decoder_decoded_T_57};
  wire [19:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_8 = {id_ctrl_decoder_decoded_orMatrixOutputs_hi_2,
    id_ctrl_decoder_decoded_orMatrixOutputs_lo_1};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_9 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_8;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_10 = |_id_ctrl_decoder_decoded_T_123;
  wire [7:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_11 = {_id_ctrl_decoder_decoded_T_25,
    _id_ctrl_decoder_decoded_T_29,_id_ctrl_decoder_decoded_T_65,_id_ctrl_decoder_decoded_T_157,
    _id_ctrl_decoder_decoded_T_159,_id_ctrl_decoder_decoded_T_169,_id_ctrl_decoder_decoded_T_185,
    _id_ctrl_decoder_decoded_T_191};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_12 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_11;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_13 = |_id_ctrl_decoder_decoded_T_25;
  wire [6:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_14 = {_id_ctrl_decoder_decoded_T_25,
    _id_ctrl_decoder_decoded_T_29,_id_ctrl_decoder_decoded_T_73,_id_ctrl_decoder_decoded_T_153,
    _id_ctrl_decoder_decoded_T_155,_id_ctrl_decoder_decoded_T_157,_id_ctrl_decoder_decoded_T_169};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_15 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_14;
  wire [7:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_16 = {_id_ctrl_decoder_decoded_T_25,
    _id_ctrl_decoder_decoded_T_29,_id_ctrl_decoder_decoded_T_153,_id_ctrl_decoder_decoded_T_155,
    _id_ctrl_decoder_decoded_T_157,_id_ctrl_decoder_decoded_T_169,_id_ctrl_decoder_decoded_T_183,
    _id_ctrl_decoder_decoded_T_189};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_17 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_16;
  wire [4:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_18 = {_id_ctrl_decoder_decoded_T_19,
    _id_ctrl_decoder_decoded_T_45,_id_ctrl_decoder_decoded_T_71,_id_ctrl_decoder_decoded_T_151,
    _id_ctrl_decoder_decoded_T_161};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_19 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_18;
  wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_20 = {_id_ctrl_decoder_decoded_T_131,
    _id_ctrl_decoder_decoded_T_151,_id_ctrl_decoder_decoded_T_165};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_21 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_20;
  wire [4:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_22 = {_id_ctrl_decoder_decoded_T_45,
    _id_ctrl_decoder_decoded_T_129,_id_ctrl_decoder_decoded_T_131,_id_ctrl_decoder_decoded_T_143,
    _id_ctrl_decoder_decoded_T_175};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_23 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_22;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_24 = |_id_ctrl_decoder_decoded_T_75;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_25 = |_id_ctrl_decoder_decoded_T_143;
  wire [7:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_26 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_7,
    _id_ctrl_decoder_decoded_T_45,_id_ctrl_decoder_decoded_T_59,_id_ctrl_decoder_decoded_T_75,
    _id_ctrl_decoder_decoded_T_129,_id_ctrl_decoder_decoded_T_133,_id_ctrl_decoder_decoded_T_149};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_27 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_26;
  wire [6:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_28 = {_id_ctrl_decoder_decoded_T_47,
    _id_ctrl_decoder_decoded_T_53,_id_ctrl_decoder_decoded_T_95,_id_ctrl_decoder_decoded_T_103,
    _id_ctrl_decoder_decoded_T_107,_id_ctrl_decoder_decoded_T_121,_id_ctrl_decoder_decoded_T_125};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_29 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_28;
  wire [8:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_30 = {_id_ctrl_decoder_decoded_T_33,
    _id_ctrl_decoder_decoded_T_85,_id_ctrl_decoder_decoded_T_87,_id_ctrl_decoder_decoded_T_111,
    _id_ctrl_decoder_decoded_T_113,_id_ctrl_decoder_decoded_T_117,_id_ctrl_decoder_decoded_T_127,
    _id_ctrl_decoder_decoded_T_163,_id_ctrl_decoder_decoded_T_167};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_31 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_30;
  wire [5:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_32 = {_id_ctrl_decoder_decoded_T_67,
    _id_ctrl_decoder_decoded_T_77,_id_ctrl_decoder_decoded_T_89,_id_ctrl_decoder_decoded_T_91,
    _id_ctrl_decoder_decoded_T_93,_id_ctrl_decoder_decoded_T_99};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_33 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_32;
  wire [4:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_34 = {_id_ctrl_decoder_decoded_T_69,
    _id_ctrl_decoder_decoded_T_79,_id_ctrl_decoder_decoded_T_93,_id_ctrl_decoder_decoded_T_163,
    _id_ctrl_decoder_decoded_T_167};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_35 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_34;
  wire [8:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_12 = {_id_ctrl_decoder_decoded_T_57,
    _id_ctrl_decoder_decoded_T_59,_id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_75,
    _id_ctrl_decoder_decoded_T_81,_id_ctrl_decoder_decoded_T_95,_id_ctrl_decoder_decoded_T_129,
    _id_ctrl_decoder_decoded_T_131,_id_ctrl_decoder_decoded_T_143};
  wire [17:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_36 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_3
    ,_id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_11,_id_ctrl_decoder_decoded_T_21,
    _id_ctrl_decoder_decoded_T_23,_id_ctrl_decoder_decoded_T_37,_id_ctrl_decoder_decoded_T_39,
    _id_ctrl_decoder_decoded_T_47,id_ctrl_decoder_decoded_orMatrixOutputs_lo_12};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_37 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_36;
  wire [3:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_38 = {_id_ctrl_decoder_decoded_T_31,
    _id_ctrl_decoder_decoded_T_39,_id_ctrl_decoder_decoded_T_105,_id_ctrl_decoder_decoded_T_115};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_39 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_38;
  wire [1:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_40 = {_id_ctrl_decoder_decoded_T_11,
    _id_ctrl_decoder_decoded_T_39};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_41 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_40;
  wire [8:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_42 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_3,
    _id_ctrl_decoder_decoded_T_37,_id_ctrl_decoder_decoded_T_49,_id_ctrl_decoder_decoded_T_61,
    _id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_97,_id_ctrl_decoder_decoded_T_109,
    _id_ctrl_decoder_decoded_T_119};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_43 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_42;
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_17 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_3,
    _id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_21,_id_ctrl_decoder_decoded_T_23,
    _id_ctrl_decoder_decoded_T_35,_id_ctrl_decoder_decoded_T_47,_id_ctrl_decoder_decoded_T_55,
    _id_ctrl_decoder_decoded_T_59,_id_ctrl_decoder_decoded_T_67};
  wire [18:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_44 = {id_ctrl_decoder_decoded_orMatrixOutputs_hi_17,
    _id_ctrl_decoder_decoded_T_75,_id_ctrl_decoder_decoded_T_83,_id_ctrl_decoder_decoded_T_93,
    _id_ctrl_decoder_decoded_T_95,_id_ctrl_decoder_decoded_T_129,_id_ctrl_decoder_decoded_T_131,
    _id_ctrl_decoder_decoded_T_145,_id_ctrl_decoder_decoded_T_185,_id_ctrl_decoder_decoded_T_191};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_45 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_44;
  wire [1:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_46 = {_id_ctrl_decoder_decoded_T_13,
    _id_ctrl_decoder_decoded_T_39};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_47 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_46;
  wire [5:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_16 = {_id_ctrl_decoder_decoded_T_49,
    _id_ctrl_decoder_decoded_T_59,_id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_97,
    _id_ctrl_decoder_decoded_T_109,_id_ctrl_decoder_decoded_T_119};
  wire [11:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_48 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_3
    ,_id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_11,_id_ctrl_decoder_decoded_T_37,
    _id_ctrl_decoder_decoded_T_39,id_ctrl_decoder_decoded_orMatrixOutputs_lo_16};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_49 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_48;
  wire [6:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_17 = {_id_ctrl_decoder_decoded_T_35,
    _id_ctrl_decoder_decoded_T_47,_id_ctrl_decoder_decoded_T_59,_id_ctrl_decoder_decoded_T_67,
    _id_ctrl_decoder_decoded_T_95,_id_ctrl_decoder_decoded_T_105,_id_ctrl_decoder_decoded_T_115};
  wire [13:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_50 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_3
    ,_id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_11,_id_ctrl_decoder_decoded_T_21,
    _id_ctrl_decoder_decoded_T_23,_id_ctrl_decoder_decoded_T_31,id_ctrl_decoder_decoded_orMatrixOutputs_lo_17};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_51 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_50;
  wire [9:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_54 = {_id_ctrl_decoder_decoded_T_15,
    _id_ctrl_decoder_decoded_T_17,_id_ctrl_decoder_decoded_T_21,_id_ctrl_decoder_decoded_T_23,
    _id_ctrl_decoder_decoded_T_75,_id_ctrl_decoder_decoded_T_93,_id_ctrl_decoder_decoded_T_101,
    _id_ctrl_decoder_decoded_T_129,_id_ctrl_decoder_decoded_T_131,_id_ctrl_decoder_decoded_T_147};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_55 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_54;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_56 = |_id_ctrl_decoder_decoded_T_37;
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_57 = |_id_ctrl_decoder_decoded_T_39;
  wire [1:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_58 = {_id_ctrl_decoder_decoded_T_31,
    _id_ctrl_decoder_decoded_T_93};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_59 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_58;
  wire [9:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_60 = {_id_ctrl_decoder_decoded_T_25,
    _id_ctrl_decoder_decoded_T_29,_id_ctrl_decoder_decoded_T_63,_id_ctrl_decoder_decoded_T_153,
    _id_ctrl_decoder_decoded_T_155,_id_ctrl_decoder_decoded_T_157,_id_ctrl_decoder_decoded_T_169,
    _id_ctrl_decoder_decoded_T_181,_id_ctrl_decoder_decoded_T_187,_id_ctrl_decoder_decoded_T_189};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_61 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_60;
  wire [7:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_13 = {_id_ctrl_decoder_decoded_T_153,
    _id_ctrl_decoder_decoded_T_155,_id_ctrl_decoder_decoded_T_157,_id_ctrl_decoder_decoded_T_169,
    _id_ctrl_decoder_decoded_T_173,_id_ctrl_decoder_decoded_T_181,_id_ctrl_decoder_decoded_T_187,
    _id_ctrl_decoder_decoded_T_189};
  wire [7:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_16 = {_id_ctrl_decoder_decoded_T_35,
    _id_ctrl_decoder_decoded_T_39,_id_ctrl_decoder_decoded_T_43,_id_ctrl_decoder_decoded_T_47,
    _id_ctrl_decoder_decoded_T_51,_id_ctrl_decoder_decoded_T_59,_id_ctrl_decoder_decoded_T_67,
    _id_ctrl_decoder_decoded_T_75};
  wire [16:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_23 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_3
    ,_id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_9,_id_ctrl_decoder_decoded_T_11,
    _id_ctrl_decoder_decoded_T_21,_id_ctrl_decoder_decoded_T_23,_id_ctrl_decoder_decoded_T_27,
    _id_ctrl_decoder_decoded_T_29,id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_16};
  wire [32:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_62 = {id_ctrl_decoder_decoded_orMatrixOutputs_hi_23,
    _id_ctrl_decoder_decoded_T_81,_id_ctrl_decoder_decoded_T_93,_id_ctrl_decoder_decoded_T_95,
    _id_ctrl_decoder_decoded_T_129,_id_ctrl_decoder_decoded_T_133,_id_ctrl_decoder_decoded_T_137,
    _id_ctrl_decoder_decoded_T_141,_id_ctrl_decoder_decoded_T_149,id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_13};
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_63 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_62;
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_14 = {1'h0,_id_ctrl_decoder_decoded_orMatrixOutputs_T_10,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_9,_id_ctrl_decoder_decoded_orMatrixOutputs_T_7,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_5,_id_ctrl_decoder_decoded_orMatrixOutputs_T_4,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_3,_id_ctrl_decoder_decoded_orMatrixOutputs_T_2,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_1,1'h0};
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_18 = {_id_ctrl_decoder_decoded_orMatrixOutputs_T_27,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_25,_id_ctrl_decoder_decoded_orMatrixOutputs_T_24,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_23,_id_ctrl_decoder_decoded_orMatrixOutputs_T_21,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_19,_id_ctrl_decoder_decoded_orMatrixOutputs_T_17,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_15,_id_ctrl_decoder_decoded_orMatrixOutputs_T_13,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_12};
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_17 = {_id_ctrl_decoder_decoded_orMatrixOutputs_T_47,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_45,_id_ctrl_decoder_decoded_orMatrixOutputs_T_43,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_41,_id_ctrl_decoder_decoded_orMatrixOutputs_T_39,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_37,_id_ctrl_decoder_decoded_orMatrixOutputs_T_35,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_33,_id_ctrl_decoder_decoded_orMatrixOutputs_T_31,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_29};
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6 = {_id_ctrl_decoder_decoded_orMatrixOutputs_T_55,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_45,1'h0,_id_ctrl_decoder_decoded_orMatrixOutputs_T_51,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_49};
  wire [40:0] id_ctrl_decoder_decoded_orMatrixOutputs = {_id_ctrl_decoder_decoded_orMatrixOutputs_T_63,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_61,1'h0,_id_ctrl_decoder_decoded_orMatrixOutputs_T_59,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_57,_id_ctrl_decoder_decoded_orMatrixOutputs_T_56,
    id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6,id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_17,
    id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_18,id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_14};
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[9],
    id_ctrl_decoder_decoded_orMatrixOutputs[8],id_ctrl_decoder_decoded_orMatrixOutputs[7],
    id_ctrl_decoder_decoded_orMatrixOutputs[6],id_ctrl_decoder_decoded_orMatrixOutputs[5],
    id_ctrl_decoder_decoded_orMatrixOutputs[4],id_ctrl_decoder_decoded_orMatrixOutputs[3],
    id_ctrl_decoder_decoded_orMatrixOutputs[2],id_ctrl_decoder_decoded_orMatrixOutputs[1],
    id_ctrl_decoder_decoded_orMatrixOutputs[0]};
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi = {id_ctrl_decoder_decoded_orMatrixOutputs[19],
    id_ctrl_decoder_decoded_orMatrixOutputs[18],id_ctrl_decoder_decoded_orMatrixOutputs[17],
    id_ctrl_decoder_decoded_orMatrixOutputs[16],id_ctrl_decoder_decoded_orMatrixOutputs[15],
    id_ctrl_decoder_decoded_orMatrixOutputs[14],id_ctrl_decoder_decoded_orMatrixOutputs[13],
    id_ctrl_decoder_decoded_orMatrixOutputs[12],id_ctrl_decoder_decoded_orMatrixOutputs[11],
    id_ctrl_decoder_decoded_orMatrixOutputs[10]};
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[29],
    id_ctrl_decoder_decoded_orMatrixOutputs[28],id_ctrl_decoder_decoded_orMatrixOutputs[27],
    id_ctrl_decoder_decoded_orMatrixOutputs[26],id_ctrl_decoder_decoded_orMatrixOutputs[25],
    id_ctrl_decoder_decoded_orMatrixOutputs[24],id_ctrl_decoder_decoded_orMatrixOutputs[23],
    id_ctrl_decoder_decoded_orMatrixOutputs[22],id_ctrl_decoder_decoded_orMatrixOutputs[21],
    id_ctrl_decoder_decoded_orMatrixOutputs[20]};
  wire [4:0] id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[34],
    id_ctrl_decoder_decoded_orMatrixOutputs[33],id_ctrl_decoder_decoded_orMatrixOutputs[32],
    id_ctrl_decoder_decoded_orMatrixOutputs[31],id_ctrl_decoder_decoded_orMatrixOutputs[30]};
  wire [40:0] id_ctrl_decoder_decoded_invMatrixOutputs = {id_ctrl_decoder_decoded_orMatrixOutputs[40],
    id_ctrl_decoder_decoded_orMatrixOutputs[39],id_ctrl_decoder_decoded_orMatrixOutputs[38],
    id_ctrl_decoder_decoded_orMatrixOutputs[37],id_ctrl_decoder_decoded_orMatrixOutputs[36],
    id_ctrl_decoder_decoded_orMatrixOutputs[35],id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo,
    id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo,id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi,
    id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo};
  wire  id_ctrl_decoder_0 = id_ctrl_decoder_decoded_invMatrixOutputs[40];
  wire  id_ctrl_decoder_1 = id_ctrl_decoder_decoded_invMatrixOutputs[39];
  wire  id_ctrl_decoder_2 = id_ctrl_decoder_decoded_invMatrixOutputs[38];
  wire  id_ctrl_decoder_3 = id_ctrl_decoder_decoded_invMatrixOutputs[37];
  wire  id_ctrl_decoder_4 = id_ctrl_decoder_decoded_invMatrixOutputs[36];
  wire  id_ctrl_decoder_5 = id_ctrl_decoder_decoded_invMatrixOutputs[35];
  wire  id_ctrl_decoder_6 = id_ctrl_decoder_decoded_invMatrixOutputs[34];
  wire  id_ctrl_decoder_7 = id_ctrl_decoder_decoded_invMatrixOutputs[33];
  wire  id_ctrl_decoder_8 = id_ctrl_decoder_decoded_invMatrixOutputs[32];
  wire [1:0] id_ctrl_decoder_9 = id_ctrl_decoder_decoded_invMatrixOutputs[31:30];
  wire [1:0] id_ctrl_decoder_10 = id_ctrl_decoder_decoded_invMatrixOutputs[29:28];
  wire [2:0] id_ctrl_decoder_11 = id_ctrl_decoder_decoded_invMatrixOutputs[27:25];
  wire [3:0] id_ctrl_decoder_13 = id_ctrl_decoder_decoded_invMatrixOutputs[23:20];
  wire  id_ctrl_decoder_14 = id_ctrl_decoder_decoded_invMatrixOutputs[19];
  wire [4:0] id_ctrl_decoder_15 = id_ctrl_decoder_decoded_invMatrixOutputs[18:14];
  wire  id_ctrl_decoder_16 = id_ctrl_decoder_decoded_invMatrixOutputs[13];
  wire  id_ctrl_decoder_17 = id_ctrl_decoder_decoded_invMatrixOutputs[12];
  wire  id_ctrl_decoder_19 = id_ctrl_decoder_decoded_invMatrixOutputs[10];
  wire  id_ctrl_decoder_20 = id_ctrl_decoder_decoded_invMatrixOutputs[9];
  wire  id_ctrl_decoder_21 = id_ctrl_decoder_decoded_invMatrixOutputs[8];
  wire  id_ctrl_decoder_22 = id_ctrl_decoder_decoded_invMatrixOutputs[7];
  wire [2:0] id_ctrl_decoder_23 = id_ctrl_decoder_decoded_invMatrixOutputs[6:4];
  wire  id_ctrl_decoder_24 = id_ctrl_decoder_decoded_invMatrixOutputs[3];
  wire  id_ctrl_decoder_25 = id_ctrl_decoder_decoded_invMatrixOutputs[2];
  wire  id_ctrl_decoder_26 = id_ctrl_decoder_decoded_invMatrixOutputs[1];
  wire  id_ctrl_decoder_27 = id_ctrl_decoder_decoded_invMatrixOutputs[0];
  wire [4:0] id_raddr3 = ibuf_io_inst_0_bits_inst_rs3;
  wire [4:0] id_raddr2 = ibuf_io_inst_0_bits_inst_rs2;
  wire [4:0] id_raddr1 = ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0] id_waddr = ibuf_io_inst_0_bits_inst_rd;
  reg  id_reg_fence;
  wire [31:0] _id_rs_T_4 = rf_id_rs_MPORT_data;
  wire [31:0] _id_rs_T_9 = rf_id_rs_MPORT_1_data;
  wire  _id_csr_en_T = id_ctrl_decoder_23 == 3'h6;
  wire  _id_csr_en_T_1 = id_ctrl_decoder_23 == 3'h7;
  wire  _id_csr_en_T_2 = id_ctrl_decoder_23 == 3'h5;
  wire  _id_csr_en_T_3 = _id_csr_en_T | _id_csr_en_T_1;
  wire  id_csr_en = _id_csr_en_T | _id_csr_en_T_1 | _id_csr_en_T_2;
  wire  id_system_insn = id_ctrl_decoder_23 == 3'h4;
  wire  id_csr_ren = _id_csr_en_T_3 & ibuf_io_inst_0_bits_inst_rs1 == 5'h0;
  wire  _id_csr_flush_T = ~id_csr_ren;
  wire  id_csr_flush = id_system_insn | id_csr_en & ~id_csr_ren & csr_io_decode_0_write_flush;
  wire  _id_illegal_insn_T_4 = (id_ctrl_decoder_20 | id_ctrl_decoder_21) & ~csr_io_status_isa[12];
  wire  _id_illegal_insn_T_5 = ~id_ctrl_decoder_0 | _id_illegal_insn_T_4;
  wire  _id_illegal_insn_T_8 = id_ctrl_decoder_26 & ~csr_io_status_isa[0];
  wire  _id_illegal_insn_T_9 = _id_illegal_insn_T_5 | _id_illegal_insn_T_8;
  wire  _id_illegal_insn_T_11 = id_ctrl_decoder_1 & (csr_io_decode_0_fp_illegal | io_fpu_illegal_rm);
  wire  _id_illegal_insn_T_12 = _id_illegal_insn_T_9 | _id_illegal_insn_T_11;
  wire  _id_illegal_insn_T_15 = id_ctrl_decoder_27 & ~csr_io_status_isa[3];
  wire  _id_illegal_insn_T_16 = _id_illegal_insn_T_12 | _id_illegal_insn_T_15;
  wire  _id_illegal_insn_T_18 = ~csr_io_status_isa[2];
  wire  _id_illegal_insn_T_19 = ibuf_io_inst_0_bits_rvc & ~csr_io_status_isa[2];
  wire  _id_illegal_insn_T_20 = _id_illegal_insn_T_16 | _id_illegal_insn_T_19;
  wire  _id_illegal_insn_T_33 = id_ctrl_decoder_2 & csr_io_decode_0_rocc_illegal;
  wire  _id_illegal_insn_T_34 = _id_illegal_insn_T_20 | _id_illegal_insn_T_33;
  wire  _id_illegal_insn_T_38 = _id_illegal_insn_T_34 | id_ctrl_decoder_8;
  wire  _id_illegal_insn_T_42 = id_csr_en & (csr_io_decode_0_read_illegal | _id_csr_flush_T &
    csr_io_decode_0_write_illegal);
  wire  _id_illegal_insn_T_43 = _id_illegal_insn_T_38 | _id_illegal_insn_T_42;
  wire  _id_illegal_insn_T_46 = ~ibuf_io_inst_0_bits_rvc & (id_system_insn & csr_io_decode_0_system_illegal);
  wire  id_illegal_insn = _id_illegal_insn_T_43 | _id_illegal_insn_T_46;
  wire  id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26];
  wire  id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25];
  wire [3:0] id_fence_succ = ibuf_io_inst_0_bits_inst_bits[23:20];
  wire  id_fence_next = id_ctrl_decoder_25 | id_ctrl_decoder_26 & id_amo_aq;
  wire  id_mem_busy = ~io_dmem_ordered | io_dmem_req_valid;
  wire  _GEN_0 = ~id_mem_busy ? 1'h0 : id_reg_fence;
  wire  id_do_fence_x9 = id_mem_busy & (id_ctrl_decoder_26 & id_amo_rl | id_ctrl_decoder_24 | id_reg_fence & (
    id_ctrl_decoder_14 | id_ctrl_decoder_2));
  wire  id_xcpt = csr_io_interrupt | bpu_io_debug_if | bpu_io_xcpt_if | ibuf_io_inst_0_bits_xcpt0_pf_inst |
    ibuf_io_inst_0_bits_xcpt0_ae_inst | ibuf_io_inst_0_bits_xcpt1_pf_inst | ibuf_io_inst_0_bits_xcpt1_gf_inst |
    ibuf_io_inst_0_bits_xcpt1_ae_inst | id_illegal_insn;
  wire [4:0] _T_11 = ibuf_io_inst_0_bits_xcpt1_ae_inst ? 5'h1 : 5'h2;
  wire [4:0] _T_12 = ibuf_io_inst_0_bits_xcpt1_gf_inst ? 5'h14 : _T_11;
  wire [4:0] _T_13 = ibuf_io_inst_0_bits_xcpt1_pf_inst ? 5'hc : _T_12;
  wire [4:0] _T_14 = ibuf_io_inst_0_bits_xcpt0_ae_inst ? 5'h1 : _T_13;
  wire [4:0] _T_16 = ibuf_io_inst_0_bits_xcpt0_pf_inst ? 5'hc : _T_14;
  wire [4:0] _T_17 = bpu_io_xcpt_if ? 5'h3 : _T_16;
  wire [4:0] _T_18 = bpu_io_debug_if ? 5'he : _T_17;
  wire [4:0] ex_waddr = ex_reg_inst[11:7];
  wire [4:0] mem_waddr = mem_reg_inst[11:7];
  wire [4:0] wb_waddr = wb_reg_inst[11:7];
  wire  _T_29 = ex_reg_valid & ex_ctrl_wxd;
  wire  _T_30 = mem_reg_valid & mem_ctrl_wxd;
  wire  _T_32 = mem_reg_valid & mem_ctrl_wxd & ~mem_ctrl_mem;
  wire  id_bypass_src_0_0 = 5'h0 == id_raddr1;
  wire  id_bypass_src_0_1 = _T_29 & ex_waddr == id_raddr1;
  wire  id_bypass_src_0_2 = _T_32 & mem_waddr == id_raddr1;
  wire  id_bypass_src_0_3 = _T_30 & mem_waddr == id_raddr1;
  wire  id_bypass_src_1_0 = 5'h0 == id_raddr2;
  wire  id_bypass_src_1_1 = _T_29 & ex_waddr == id_raddr2;
  wire  id_bypass_src_1_2 = _T_32 & mem_waddr == id_raddr2;
  wire  id_bypass_src_1_3 = _T_30 & mem_waddr == id_raddr2;
  reg  ex_reg_rs_bypass_0;
  reg  ex_reg_rs_bypass_1;
  reg [1:0] ex_reg_rs_lsb_0;
  reg [1:0] ex_reg_rs_lsb_1;
  reg [29:0] ex_reg_rs_msb_0;
  reg [29:0] ex_reg_rs_msb_1;
  wire [31:0] _ex_rs_T_1 = ex_reg_rs_lsb_0 == 2'h1 ? mem_reg_wdata : 32'h0;
  wire [31:0] _ex_rs_T_3 = ex_reg_rs_lsb_0 == 2'h2 ? wb_reg_wdata : _ex_rs_T_1;
  wire [31:0] _ex_rs_T_5 = ex_reg_rs_lsb_0 == 2'h3 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_3;
  wire [31:0] _ex_rs_T_6 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0};
  wire [31:0] _ex_rs_T_8 = ex_reg_rs_lsb_1 == 2'h1 ? mem_reg_wdata : 32'h0;
  wire [31:0] _ex_rs_T_10 = ex_reg_rs_lsb_1 == 2'h2 ? wb_reg_wdata : _ex_rs_T_8;
  wire [31:0] _ex_rs_T_12 = ex_reg_rs_lsb_1 == 2'h3 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_10;
  wire [31:0] _ex_rs_T_13 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1};
  wire [31:0] ex_rs_1 = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13;
  wire  _ex_imm_sign_T = ex_ctrl_sel_imm == 3'h5;
  wire  _ex_imm_sign_T_2 = ex_reg_inst[31];
  wire  ex_imm_sign = ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2);
  wire  _ex_imm_b30_20_T = ex_ctrl_sel_imm == 3'h2;
  wire [10:0] _ex_imm_b30_20_T_2 = ex_reg_inst[30:20];
  wire [7:0] _ex_imm_b19_12_T_4 = ex_reg_inst[19:12];
  wire  _ex_imm_b11_T_2 = _ex_imm_b30_20_T | _ex_imm_sign_T;
  wire  _ex_imm_b11_T_5 = ex_reg_inst[20];
  wire  _ex_imm_b11_T_6 = ex_ctrl_sel_imm == 3'h1;
  wire  _ex_imm_b11_T_8 = ex_reg_inst[7];
  wire  _ex_imm_b11_T_9 = ex_ctrl_sel_imm == 3'h1 ? $signed(_ex_imm_b11_T_8) : $signed(ex_imm_sign);
  wire  _ex_imm_b11_T_10 = ex_ctrl_sel_imm == 3'h3 ? $signed(_ex_imm_b11_T_5) : $signed(_ex_imm_b11_T_9);
  wire [5:0] ex_imm_b10_5 = _ex_imm_b11_T_2 ? 6'h0 : ex_reg_inst[30:25];
  wire  _ex_imm_b4_1_T_1 = ex_ctrl_sel_imm == 3'h0;
  wire [3:0] _ex_imm_b4_1_T_8 = _ex_imm_sign_T ? ex_reg_inst[19:16] : ex_reg_inst[24:21];
  wire [3:0] _ex_imm_b4_1_T_9 = ex_ctrl_sel_imm == 3'h0 | _ex_imm_b11_T_6 ? ex_reg_inst[11:8] : _ex_imm_b4_1_T_8;
  wire [3:0] ex_imm_b4_1 = _ex_imm_b30_20_T ? 4'h0 : _ex_imm_b4_1_T_9;
  wire  _ex_imm_b0_T_6 = _ex_imm_sign_T & ex_reg_inst[15];
  wire  _ex_imm_b0_T_7 = ex_ctrl_sel_imm == 3'h4 ? ex_reg_inst[20] : _ex_imm_b0_T_6;
  wire  ex_imm_b0 = _ex_imm_b4_1_T_1 ? ex_reg_inst[7] : _ex_imm_b0_T_7;
  wire  ex_imm_hi_lo_lo = _ex_imm_b30_20_T | _ex_imm_sign_T ? $signed(1'sh0) : $signed(_ex_imm_b11_T_10);
  wire [7:0] ex_imm_hi_lo_hi = ex_ctrl_sel_imm != 3'h2 & ex_ctrl_sel_imm != 3'h3 ? $signed({8{ex_imm_sign}}) : $signed(
    _ex_imm_b19_12_T_4);
  wire [10:0] ex_imm_hi_hi_lo = ex_ctrl_sel_imm == 3'h2 ? $signed(_ex_imm_b30_20_T_2) : $signed({11{ex_imm_sign}});
  wire  ex_imm_hi_hi_hi = ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2);
  wire [31:0] ex_imm = {ex_imm_hi_hi_hi,ex_imm_hi_hi_lo,ex_imm_hi_lo_hi,ex_imm_hi_lo_lo,ex_imm_b10_5,ex_imm_b4_1,
    ex_imm_b0};
  wire [31:0] _ex_op1_T = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6;
  wire [31:0] _ex_op1_T_3 = 2'h1 == ex_ctrl_sel_alu1 ? $signed(_ex_op1_T) : $signed(32'sh0);
  wire [31:0] _ex_op2_T = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13;
  wire [3:0] _ex_op2_T_1 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  wire [31:0] _ex_op2_T_3 = 2'h2 == ex_ctrl_sel_alu2 ? $signed(_ex_op2_T) : $signed(32'sh0);
  wire [31:0] _ex_op2_T_5 = 2'h3 == ex_ctrl_sel_alu2 ? $signed(ex_imm) : $signed(_ex_op2_T_3);
  wire  _T_144 = id_raddr1 != 5'h0;
  wire  _T_145 = id_ctrl_decoder_7 & id_raddr1 != 5'h0;
  wire  _data_hazard_ex_T = id_raddr1 == ex_waddr;
  wire  _T_146 = id_raddr2 != 5'h0;
  wire  _T_147 = id_ctrl_decoder_6 & id_raddr2 != 5'h0;
  wire  _data_hazard_ex_T_2 = id_raddr2 == ex_waddr;
  wire  _T_149 = id_ctrl_decoder_22 & id_waddr != 5'h0;
  wire  _data_hazard_ex_T_4 = id_waddr == ex_waddr;
  wire  _data_hazard_ex_T_7 = _T_145 & _data_hazard_ex_T | _T_147 & _data_hazard_ex_T_2 | _T_149 & _data_hazard_ex_T_4;
  wire  data_hazard_ex = ex_ctrl_wxd & _data_hazard_ex_T_7;
  wire  ex_cannot_bypass = ex_ctrl_csr != 3'h0 | ex_ctrl_jalr | ex_ctrl_mem | ex_ctrl_mul | ex_ctrl_div | ex_ctrl_fp |
    ex_ctrl_rocc;
  wire  _fp_data_hazard_ex_T_5 = id_raddr3 == ex_waddr;
  wire  _fp_data_hazard_ex_T_11 = io_fpu_dec_ren1 & _data_hazard_ex_T | io_fpu_dec_ren2 & _data_hazard_ex_T_2 |
    io_fpu_dec_ren3 & _fp_data_hazard_ex_T_5 | io_fpu_dec_wen & _data_hazard_ex_T_4;
  wire  fp_data_hazard_ex = id_ctrl_decoder_1 & ex_ctrl_wfd & _fp_data_hazard_ex_T_11;
  wire  id_ex_hazard = ex_reg_valid & (data_hazard_ex & ex_cannot_bypass | fp_data_hazard_ex);
  wire  _data_hazard_mem_T = id_raddr1 == mem_waddr;
  wire  _data_hazard_mem_T_2 = id_raddr2 == mem_waddr;
  wire  _data_hazard_mem_T_4 = id_waddr == mem_waddr;
  wire  _data_hazard_mem_T_7 = _T_145 & _data_hazard_mem_T | _T_147 & _data_hazard_mem_T_2 | _T_149 &
    _data_hazard_mem_T_4;
  wire  data_hazard_mem = mem_ctrl_wxd & _data_hazard_mem_T_7;
  wire  mem_cannot_bypass = mem_ctrl_csr != 3'h0 | mem_ctrl_mem & mem_reg_slow_bypass | mem_ctrl_mul | mem_ctrl_div |
    mem_ctrl_fp | mem_ctrl_rocc;
  wire  _fp_data_hazard_mem_T_5 = id_raddr3 == mem_waddr;
  wire  _fp_data_hazard_mem_T_11 = io_fpu_dec_ren1 & _data_hazard_mem_T | io_fpu_dec_ren2 & _data_hazard_mem_T_2 |
    io_fpu_dec_ren3 & _fp_data_hazard_mem_T_5 | io_fpu_dec_wen & _data_hazard_mem_T_4;
  wire  fp_data_hazard_mem = id_ctrl_decoder_1 & mem_ctrl_wfd & _fp_data_hazard_mem_T_11;
  wire  id_mem_hazard = mem_reg_valid & (data_hazard_mem & mem_cannot_bypass | fp_data_hazard_mem);
  wire  _data_hazard_wb_T = id_raddr1 == wb_waddr;
  wire  _data_hazard_wb_T_2 = id_raddr2 == wb_waddr;
  wire  _data_hazard_wb_T_4 = id_waddr == wb_waddr;
  wire  _data_hazard_wb_T_7 = _T_145 & _data_hazard_wb_T | _T_147 & _data_hazard_wb_T_2 | _T_149 & _data_hazard_wb_T_4;
  wire  data_hazard_wb = wb_ctrl_wxd & _data_hazard_wb_T_7;
  wire  wb_dcache_miss = wb_ctrl_mem & ~io_dmem_resp_valid;
  wire  wb_set_sboard = wb_ctrl_div | wb_dcache_miss | wb_ctrl_rocc;
  wire  _fp_data_hazard_wb_T_5 = id_raddr3 == wb_waddr;
  wire  _fp_data_hazard_wb_T_11 = io_fpu_dec_ren1 & _data_hazard_wb_T | io_fpu_dec_ren2 & _data_hazard_wb_T_2 |
    io_fpu_dec_ren3 & _fp_data_hazard_wb_T_5 | io_fpu_dec_wen & _data_hazard_wb_T_4;
  wire  fp_data_hazard_wb = id_ctrl_decoder_1 & wb_ctrl_wfd & _fp_data_hazard_wb_T_11;
  wire  id_wb_hazard = wb_reg_valid & (data_hazard_wb & wb_set_sboard | fp_data_hazard_wb);
  reg [31:0] _r;
  wire [31:0] r = {_r[31:1], 1'h0};
  wire [31:0] _id_sboard_hazard_T = r >> id_raddr1;
  wire  dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  wire  dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
  wire  dmem_resp_xpu = ~io_dmem_resp_bits_tag[0];
  wire  ll_wen_x2 = div_io_resp_ready & div_io_resp_valid;
  wire  ll_wen = dmem_resp_replay & dmem_resp_xpu | ll_wen_x2;
  wire [4:0] dmem_resp_waddr = io_dmem_resp_bits_tag[5:1];
  wire [4:0] ll_waddr = dmem_resp_replay & dmem_resp_xpu ? dmem_resp_waddr : div_io_resp_bits_tag;
  wire  _id_sboard_hazard_T_3 = ll_wen & ll_waddr == id_raddr1;
  wire  _id_sboard_hazard_T_5 = _id_sboard_hazard_T[0] & ~_id_sboard_hazard_T_3;
  wire [31:0] _id_sboard_hazard_T_7 = r >> id_raddr2;
  wire  _id_sboard_hazard_T_10 = ll_wen & ll_waddr == id_raddr2;
  wire  _id_sboard_hazard_T_12 = _id_sboard_hazard_T_7[0] & ~_id_sboard_hazard_T_10;
  wire [31:0] _id_sboard_hazard_T_14 = r >> id_waddr;
  wire  _id_sboard_hazard_T_17 = ll_wen & ll_waddr == id_waddr;
  wire  _id_sboard_hazard_T_19 = _id_sboard_hazard_T_14[0] & ~_id_sboard_hazard_T_17;
  wire  id_sboard_hazard = _T_145 & _id_sboard_hazard_T_5 | _T_147 & _id_sboard_hazard_T_12 | _T_149 &
    _id_sboard_hazard_T_19;
  wire  _ctrl_stalld_T_5 = csr_io_singleStep & (ex_reg_valid | mem_reg_valid | wb_reg_valid);
  wire  _ctrl_stalld_T_6 = id_ex_hazard | id_mem_hazard | id_wb_hazard | id_sboard_hazard | _ctrl_stalld_T_5;
  wire  _ctrl_stalld_T_9 = id_csr_en & csr_io_decode_0_fp_csr & ~io_fpu_fcsr_rdy;
  wire  _ctrl_stalld_T_10 = _ctrl_stalld_T_6 | _ctrl_stalld_T_9;
  reg [31:0] id_stall_fpu__r;
  wire [31:0] _id_stall_fpu_T_18 = id_stall_fpu__r >> id_raddr1;
  wire [31:0] _id_stall_fpu_T_21 = id_stall_fpu__r >> id_raddr2;
  wire [31:0] _id_stall_fpu_T_24 = id_stall_fpu__r >> id_raddr3;
  wire [31:0] _id_stall_fpu_T_27 = id_stall_fpu__r >> id_waddr;
  wire  id_stall_fpu = io_fpu_dec_ren1 & _id_stall_fpu_T_18[0] | io_fpu_dec_ren2 & _id_stall_fpu_T_21[0] |
    io_fpu_dec_ren3 & _id_stall_fpu_T_24[0] | io_fpu_dec_wen & _id_stall_fpu_T_27[0];
  wire  _ctrl_stalld_T_11 = id_ctrl_decoder_1 & id_stall_fpu;
  wire  _ctrl_stalld_T_12 = _ctrl_stalld_T_10 | _ctrl_stalld_T_11;
  reg  blocked;
  wire  _dcache_blocked_T = ~io_dmem_perf_grant;
  wire  dcache_blocked = blocked & ~io_dmem_perf_grant;
  wire  _ctrl_stalld_T_13 = id_ctrl_decoder_14 & dcache_blocked;
  wire  _ctrl_stalld_T_14 = _ctrl_stalld_T_12 | _ctrl_stalld_T_13;
  reg  rocc_blocked;
  wire  _ctrl_stalld_T_15 = id_ctrl_decoder_2 & rocc_blocked;
  wire  _ctrl_stalld_T_16 = _ctrl_stalld_T_14 | _ctrl_stalld_T_15;
  wire  wb_wxd = wb_reg_valid & wb_ctrl_wxd;
  wire  _ctrl_stalld_T_17 = ~wb_wxd;
  wire  _ctrl_stalld_T_22 = id_ctrl_decoder_21 & (~(div_io_req_ready | div_io_resp_valid & ~wb_wxd) | div_io_req_valid);
  wire  _ctrl_stalld_T_23 = _ctrl_stalld_T_16 | _ctrl_stalld_T_22;
  wire  _ctrl_stalld_T_26 = _ctrl_stalld_T_23 | id_do_fence_x9;
  wire  _ctrl_stalld_T_27 = _ctrl_stalld_T_26 | csr_io_csr_stall;
  wire  ctrl_stalld = _ctrl_stalld_T_27 | id_reg_pause;
  wire  ctrl_killd = ~ibuf_io_inst_0_valid | ibuf_io_inst_0_bits_replay | take_pc_mem_wb | ctrl_stalld |
    csr_io_interrupt;
  wire  _ex_reg_valid_T = ~ctrl_killd;
  wire  _ex_reg_replay_T = ~take_pc_mem_wb;
  wire  _ex_reg_replay_T_1 = ~take_pc_mem_wb & ibuf_io_inst_0_valid;
  wire  _GEN_1 = id_ctrl_decoder_25 & id_fence_succ == 4'h0 | id_reg_pause;
  wire  _GEN_2 = id_fence_next | _GEN_0;
  wire [2:0] _T_37 = {ibuf_io_inst_0_bits_xcpt1_pf_inst,ibuf_io_inst_0_bits_xcpt1_gf_inst,
    ibuf_io_inst_0_bits_xcpt1_ae_inst};
  wire  _GEN_5 = |_T_37 | ibuf_io_inst_0_bits_rvc;
  wire [2:0] _T_39 = {ibuf_io_inst_0_bits_xcpt0_pf_inst,1'h0,ibuf_io_inst_0_bits_xcpt0_ae_inst};
  wire  _T_42 = id_ctrl_decoder_15 == 5'h14;
  wire  _T_43 = id_ctrl_decoder_15 == 5'h15;
  wire  _T_44 = id_ctrl_decoder_15 == 5'h16;
  wire  _T_45 = id_ctrl_decoder_15 == 5'h5;
  wire  _T_48 = _T_42 | _T_43 | _T_44 | _T_45;
  wire [1:0] _ex_reg_mem_size_T_6 = {_T_146,_T_144};
  wire  do_bypass = id_bypass_src_0_0 | id_bypass_src_0_1 | id_bypass_src_0_2 | id_bypass_src_0_3;
  wire [1:0] _bypass_src_T = id_bypass_src_0_2 ? 2'h2 : 2'h3;
  wire [1:0] _bypass_src_T_1 = id_bypass_src_0_1 ? 2'h1 : _bypass_src_T;
  wire  _wb_valid_T_2 = ~wb_xcpt;
  wire  wb_valid = wb_reg_valid & ~replay_wb & ~wb_xcpt;
  wire  wb_wen = wb_valid & wb_ctrl_wxd;
  wire  rf_wen = wb_wen | ll_wen;
  wire [4:0] rf_waddr = ll_wen ? ll_waddr : wb_waddr;
  wire  _T_139 = rf_waddr != 5'h0;
  wire  _rf_wdata_T = dmem_resp_valid & dmem_resp_xpu;
  wire [31:0] ll_wdata = div_io_resp_bits_data;
  wire [31:0] _rf_wdata_T_4 = wb_ctrl_csr != 3'h0 ? csr_io_rw_rdata : wb_reg_wdata;
  wire [31:0] _rf_wdata_T_5 = ll_wen ? ll_wdata : _rf_wdata_T_4;
  wire [31:0] rf_wdata = dmem_resp_valid & dmem_resp_xpu ? io_dmem_resp_bits_data : _rf_wdata_T_5;
  wire [31:0] _GEN_234 = rf_waddr == id_raddr1 ? rf_wdata : _id_rs_T_4;
  wire [31:0] _GEN_241 = rf_waddr != 5'h0 ? _GEN_234 : _id_rs_T_4;
  wire [31:0] id_rs_0 = rf_wen ? _GEN_241 : _id_rs_T_4;
  wire  do_bypass_1 = id_bypass_src_1_0 | id_bypass_src_1_1 | id_bypass_src_1_2 | id_bypass_src_1_3;
  wire [1:0] _bypass_src_T_2 = id_bypass_src_1_2 ? 2'h2 : 2'h3;
  wire [31:0] _GEN_235 = rf_waddr == id_raddr2 ? rf_wdata : _id_rs_T_9;
  wire [31:0] _GEN_242 = rf_waddr != 5'h0 ? _GEN_235 : _id_rs_T_9;
  wire [31:0] id_rs_1 = rf_wen ? _GEN_242 : _id_rs_T_9;
  wire [31:0] inst = ibuf_io_inst_0_bits_rvc ? {{16'd0}, ibuf_io_inst_0_bits_raw[15:0]} : ibuf_io_inst_0_bits_raw;
  wire  id_load_use = mem_reg_valid & data_hazard_mem & mem_ctrl_mem;
  wire  _replay_ex_structural_T = ~io_dmem_req_ready;
  wire  _replay_ex_structural_T_3 = ex_ctrl_div & ~div_io_req_ready;
  wire  replay_ex_structural = ex_ctrl_mem & ~io_dmem_req_ready | _replay_ex_structural_T_3;
  wire  replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  wire  replay_ex = ex_reg_replay | ex_reg_valid & (replay_ex_structural | replay_ex_load_use);
  wire  ctrl_killx = take_pc_mem_wb | replay_ex | ~ex_reg_valid;
  wire  _ex_slow_bypass_T = ex_ctrl_mem_cmd == 5'h7;
  wire  ex_slow_bypass = ex_ctrl_mem_cmd == 5'h7 | ex_reg_mem_size < 2'h2;
  wire  ex_sfence = ex_ctrl_mem & (ex_ctrl_mem_cmd == 5'h14 | ex_ctrl_mem_cmd == 5'h15 | ex_ctrl_mem_cmd == 5'h16);
  wire  ex_xcpt = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  wire  mem_pc_valid = mem_reg_valid | mem_reg_replay | mem_reg_xcpt_interrupt;
  wire  mem_npc_misaligned = _id_illegal_insn_T_18 & mem_npc[1] & ~mem_reg_sfence;
  wire [31:0] mem_int_wdata = _take_pc_mem_T & (mem_ctrl_jalr ^ mem_npc_misaligned) ? $signed(mem_br_target) : $signed(
    mem_reg_wdata);
  wire  mem_cfi = mem_ctrl_branch | mem_ctrl_jalr | mem_ctrl_jal;
  wire  mem_cfi_taken = _mem_br_target_T_1 | mem_ctrl_jalr | mem_ctrl_jal;
  wire  _mem_reg_valid_T = ~ctrl_killx;
  wire  _mem_reg_load_T = ex_ctrl_mem_cmd == 5'h0;
  wire  _mem_reg_load_T_1 = ex_ctrl_mem_cmd == 5'h10;
  wire  _mem_reg_load_T_2 = ex_ctrl_mem_cmd == 5'h6;
  wire  _mem_reg_load_T_6 = _mem_reg_load_T | _mem_reg_load_T_1 | _mem_reg_load_T_2 | _ex_slow_bypass_T;
  wire  _mem_reg_load_T_7 = ex_ctrl_mem_cmd == 5'h4;
  wire  _mem_reg_load_T_8 = ex_ctrl_mem_cmd == 5'h9;
  wire  _mem_reg_load_T_9 = ex_ctrl_mem_cmd == 5'ha;
  wire  _mem_reg_load_T_10 = ex_ctrl_mem_cmd == 5'hb;
  wire  _mem_reg_load_T_13 = _mem_reg_load_T_7 | _mem_reg_load_T_8 | _mem_reg_load_T_9 | _mem_reg_load_T_10;
  wire  _mem_reg_load_T_14 = ex_ctrl_mem_cmd == 5'h8;
  wire  _mem_reg_load_T_15 = ex_ctrl_mem_cmd == 5'hc;
  wire  _mem_reg_load_T_16 = ex_ctrl_mem_cmd == 5'hd;
  wire  _mem_reg_load_T_17 = ex_ctrl_mem_cmd == 5'he;
  wire  _mem_reg_load_T_18 = ex_ctrl_mem_cmd == 5'hf;
  wire  _mem_reg_load_T_22 = _mem_reg_load_T_14 | _mem_reg_load_T_15 | _mem_reg_load_T_16 | _mem_reg_load_T_17 |
    _mem_reg_load_T_18;
  wire  _mem_reg_load_T_23 = _mem_reg_load_T_13 | _mem_reg_load_T_22;
  wire  _mem_reg_load_T_24 = _mem_reg_load_T_6 | _mem_reg_load_T_23;
  wire  _mem_reg_store_T_22 = ex_ctrl_mem_cmd == 5'h1 | ex_ctrl_mem_cmd == 5'h11 | _ex_slow_bypass_T |
    _mem_reg_load_T_23;
  wire [31:0] _mem_reg_wdata_T = alu_io_out;
  wire [1:0] size = ex_ctrl_rocc ? 2'h2 : ex_reg_mem_size;
  wire [31:0] _mem_reg_rs2_T_3 = {ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0]};
  wire [31:0] _mem_reg_rs2_T_6 = {ex_rs_1[15:0],ex_rs_1[15:0]};
  wire [31:0] _mem_reg_rs2_T_7 = size == 2'h1 ? _mem_reg_rs2_T_6 : ex_rs_1;
  wire  _GEN_80 = ex_ctrl_jalr & csr_io_status_debug | ex_ctrl_fence_i;
  wire  _GEN_81 = ex_ctrl_jalr & csr_io_status_debug | ex_reg_flush_pipe;
  wire  mem_breakpoint = mem_reg_load & bpu_io_xcpt_ld | mem_reg_store & bpu_io_xcpt_st;
  wire  mem_debug_breakpoint = mem_reg_load & bpu_io_debug_ld | mem_reg_store & bpu_io_debug_st;
  wire  mem_ldst_xcpt = mem_debug_breakpoint | mem_breakpoint;
  wire [3:0] mem_ldst_cause = mem_debug_breakpoint ? 4'he : 4'h3;
  wire  _T_74 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  wire  _T_75 = mem_reg_valid & mem_npc_misaligned;
  wire  _T_76 = mem_reg_valid & mem_ldst_xcpt;
  wire  mem_xcpt = _T_74 | _T_75 | _T_76;
  wire [3:0] _T_78 = _T_75 ? 4'h0 : mem_ldst_cause;
  wire  dcache_kill_mem = _T_30 & io_dmem_replay_next;
  wire  fpu_kill_mem = mem_reg_valid & mem_ctrl_fp & io_fpu_nack_mem;
  wire  replay_mem = dcache_kill_mem | mem_reg_replay | fpu_kill_mem;
  wire  killm_common = dcache_kill_mem | take_pc_wb | mem_reg_xcpt | ~mem_reg_valid;
  reg  div_io_kill_REG;
  wire  ctrl_killm = killm_common | mem_xcpt | fpu_kill_mem;
  wire  _wb_reg_valid_T = ~ctrl_killm;
  wire  _wb_reg_replay_T = ~take_pc_wb;
  wire [2:0] _T_119 = _T_109 ? 3'h6 : 3'h4;
  wire [2:0] _T_120 = _T_107 ? 3'h5 : _T_119;
  wire [2:0] _T_121 = _T_105 ? 3'h7 : _T_120;
  wire [4:0] _T_122 = {{2'd0}, _T_121};
  wire [4:0] _T_124 = _T_99 ? 5'hd : _T_122;
  wire [4:0] _T_125 = _T_97 ? 5'hf : _T_124;
  wire [15:0] _csr_io_inst_0_T_3 = &wb_reg_raw_inst[1:0] ? wb_reg_inst[31:16] : 16'h0;
  wire [31:0] _io_fpu_time_T = csr_io_time;
  wire  tval_dmem_addr = ~wb_reg_xcpt;
  wire  _tval_any_addr_T = wb_reg_cause == 32'h3;
  wire  _tval_any_addr_T_1 = wb_reg_cause == 32'h1;
  wire  _tval_any_addr_T_2 = wb_reg_cause == 32'hc;
  wire  _tval_any_addr_T_3 = wb_reg_cause == 32'h14;
  wire  _tval_any_addr_T_6 = _tval_any_addr_T | _tval_any_addr_T_1 | _tval_any_addr_T_2 | _tval_any_addr_T_3;
  wire  tval_any_addr = tval_dmem_addr | _tval_any_addr_T_6;
  wire  tval_inst = wb_reg_cause == 32'h2;
  wire  tval_valid = wb_xcpt & (tval_any_addr | tval_inst);
  wire  htval_valid_imem = wb_reg_xcpt & _tval_any_addr_T_3;
  wire  _csr_io_htval_T_3 = ~reset;
  wire [2:0] _csr_io_rw_cmd_T = wb_reg_valid ? 3'h0 : 3'h4;
  wire [2:0] _csr_io_rw_cmd_T_1 = ~_csr_io_rw_cmd_T;
  wire [31:0] _T_150 = 32'h1 << ll_waddr;
  wire [31:0] _T_151 = ll_wen ? _T_150 : 32'h0;
  wire [31:0] _T_152 = ~_T_151;
  wire [31:0] _T_153 = r & _T_152;
  wire  _T_155 = wb_set_sboard & wb_wen;
  wire [31:0] _T_156 = 32'h1 << wb_waddr;
  wire [31:0] _T_157 = _T_155 ? _T_156 : 32'h0;
  wire [31:0] _T_158 = _T_153 | _T_157;
  wire  _T_159 = ll_wen | _T_155;
  wire  _id_stall_fpu_T_2 = (wb_dcache_miss & wb_ctrl_wfd | io_fpu_sboard_set) & wb_valid;
  wire [31:0] _id_stall_fpu_T_4 = _id_stall_fpu_T_2 ? _T_156 : 32'h0;
  wire [31:0] _id_stall_fpu_T_5 = id_stall_fpu__r | _id_stall_fpu_T_4;
  wire  _id_stall_fpu_T_7 = dmem_resp_replay & io_dmem_resp_bits_tag[0];
  wire [31:0] _id_stall_fpu_T_8 = 32'h1 << dmem_resp_waddr;
  wire [31:0] _id_stall_fpu_T_9 = _id_stall_fpu_T_7 ? _id_stall_fpu_T_8 : 32'h0;
  wire [31:0] _id_stall_fpu_T_10 = ~_id_stall_fpu_T_9;
  wire [31:0] _id_stall_fpu_T_11 = _id_stall_fpu_T_5 & _id_stall_fpu_T_10;
  wire  _id_stall_fpu_T_12 = _id_stall_fpu_T_2 | _id_stall_fpu_T_7;
  wire [31:0] _id_stall_fpu_T_13 = 32'h1 << io_fpu_sboard_clra;
  wire [31:0] _id_stall_fpu_T_14 = io_fpu_sboard_clr ? _id_stall_fpu_T_13 : 32'h0;
  wire [31:0] _id_stall_fpu_T_15 = ~_id_stall_fpu_T_14;
  wire [31:0] _id_stall_fpu_T_16 = _id_stall_fpu_T_11 & _id_stall_fpu_T_15;
  wire  _id_stall_fpu_T_17 = _id_stall_fpu_T_2 | _id_stall_fpu_T_7 | io_fpu_sboard_clr;
  wire [31:0] _io_imem_req_bits_pc_T_1 = replay_wb ? wb_reg_pc : mem_npc;
  wire  _io_imem_progress_T = ~replay_wb_common;
  reg  io_imem_progress_REG;
  wire  _io_imem_btb_update_bits_cfiType_T = mem_ctrl_jal | mem_ctrl_jalr;
  wire [4:0] _io_imem_btb_update_bits_cfiType_T_5 = mem_reg_inst[19:15] & 5'h1b;
  wire [1:0] _io_imem_btb_update_bits_cfiType_T_10 = mem_ctrl_jalr & 5'h1 == _io_imem_btb_update_bits_cfiType_T_5 ? 2'h3
     : {{1'd0}, _io_imem_btb_update_bits_cfiType_T};
  wire [1:0] _io_imem_btb_update_bits_br_pc_T = mem_reg_rvc ? 2'h0 : 2'h2;
  wire [31:0] _GEN_256 = {{30'd0}, _io_imem_btb_update_bits_br_pc_T};
  wire [31:0] _io_imem_btb_update_bits_pc_T = ~io_imem_btb_update_bits_br_pc;
  wire [31:0] _io_imem_btb_update_bits_pc_T_1 = _io_imem_btb_update_bits_pc_T | 32'h3;
  wire [5:0] ex_dcache_tag = {ex_waddr,ex_ctrl_fp};
  wire  unpause = csr_io_time[4:0] == 5'h0 | csr_io_inhibit_cycle | io_dmem_perf_release | take_pc_mem_wb;
  wire  coreMonitorBundle_valid = csr_io_trace_0_valid & ~csr_io_trace_0_exception;
  wire [31:0] coreMonitorBundle_pc = csr_io_trace_0_iaddr;
  wire  coreMonitorBundle_wrenx = wb_wen & ~wb_set_sboard;
  reg [31:0] coreMonitorBundle_rd0val_x23;
  reg [31:0] coreMonitorBundle_rd0val_REG;
  reg [31:0] coreMonitorBundle_rd1val_x29;
  reg [31:0] coreMonitorBundle_rd1val_REG;
  wire [4:0] _T_161 = wb_ctrl_wxd | wb_ctrl_wfd ? wb_waddr : 5'h0;
  wire [31:0] _T_162 = coreMonitorBundle_wrenx ? rf_wdata : 32'h0;
  wire  _T_163 = wb_ctrl_rxs1 | wb_ctrl_rfs1;
  wire [4:0] _T_164 = wb_ctrl_rxs1 | wb_ctrl_rfs1 ? wb_reg_inst[19:15] : 5'h0;
  wire [31:0] _T_166 = _T_163 ? coreMonitorBundle_rd0val_REG : 32'h0;
  wire  _T_167 = wb_ctrl_rxs2 | wb_ctrl_rfs2;
  wire [4:0] _T_168 = wb_ctrl_rxs2 | wb_ctrl_rfs2 ? wb_reg_inst[24:20] : 5'h0;
  wire [31:0] _T_170 = _T_167 ? coreMonitorBundle_rd1val_REG : 32'h0;
  wire [31:0] coreMonitorBundle_inst = csr_io_trace_0_insn;
  IBuf ibuf (
    .clock(ibuf_clock),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_btb_taken(ibuf_io_imem_bits_btb_taken),
    .io_imem_bits_btb_bridx(ibuf_io_imem_bits_btb_bridx),
    .io_imem_bits_btb_entry(ibuf_io_imem_bits_btb_entry),
    .io_imem_bits_btb_bht_history(ibuf_io_imem_bits_btb_bht_history),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_xcpt_pf_inst(ibuf_io_imem_bits_xcpt_pf_inst),
    .io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_btb_resp_entry(ibuf_io_btb_resp_entry),
    .io_btb_resp_bht_history(ibuf_io_btb_resp_bht_history),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_xcpt0_pf_inst(ibuf_io_inst_0_bits_xcpt0_pf_inst),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_bits_xcpt1_gf_inst(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw)
  );
  CSRFile csr (
    .clock(csr_clock),
    .reset(csr_reset),
    .io_ungated_clock(csr_io_ungated_clock),
    .io_interrupts_debug(csr_io_interrupts_debug),
    .io_interrupts_mtip(csr_io_interrupts_mtip),
    .io_interrupts_msip(csr_io_interrupts_msip),
    .io_interrupts_meip(csr_io_interrupts_meip),
    .io_interrupts_seip(csr_io_interrupts_seip),
    .io_hartid(csr_io_hartid),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_decode_0_inst(csr_io_decode_0_inst),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
    .io_decode_0_rocc_illegal(csr_io_decode_0_rocc_illegal),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_csr_stall(csr_io_csr_stall),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_cease(csr_io_status_cease),
    .io_status_wfi(csr_io_status_wfi),
    .io_status_isa(csr_io_status_isa),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_dv(csr_io_status_dv),
    .io_status_prv(csr_io_status_prv),
    .io_status_v(csr_io_status_v),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_mpv(csr_io_status_mpv),
    .io_status_gva(csr_io_status_gva),
    .io_status_mbe(csr_io_status_mbe),
    .io_status_sbe(csr_io_status_sbe),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_vs(csr_io_status_vs),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_ube(csr_io_status_ube),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_mode(csr_io_ptbr_mode),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_tval(csr_io_tval),
    .io_gva(csr_io_gva),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_action(csr_io_bp_0_control_action),
    .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_address(csr_io_bp_0_address),
    .io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
    .io_pmp_0_addr(csr_io_pmp_0_addr),
    .io_pmp_0_mask(csr_io_pmp_0_mask),
    .io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
    .io_pmp_1_addr(csr_io_pmp_1_addr),
    .io_pmp_1_mask(csr_io_pmp_1_mask),
    .io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
    .io_pmp_2_addr(csr_io_pmp_2_addr),
    .io_pmp_2_mask(csr_io_pmp_2_mask),
    .io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
    .io_pmp_3_addr(csr_io_pmp_3_addr),
    .io_pmp_3_mask(csr_io_pmp_3_mask),
    .io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
    .io_pmp_4_addr(csr_io_pmp_4_addr),
    .io_pmp_4_mask(csr_io_pmp_4_mask),
    .io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
    .io_pmp_5_addr(csr_io_pmp_5_addr),
    .io_pmp_5_mask(csr_io_pmp_5_mask),
    .io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
    .io_pmp_6_addr(csr_io_pmp_6_addr),
    .io_pmp_6_mask(csr_io_pmp_6_mask),
    .io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
    .io_pmp_7_addr(csr_io_pmp_7_addr),
    .io_pmp_7_mask(csr_io_pmp_7_mask),
    .io_inhibit_cycle(csr_io_inhibit_cycle),
    .io_inst_0(csr_io_inst_0),
    .io_trace_0_valid(csr_io_trace_0_valid),
    .io_trace_0_iaddr(csr_io_trace_0_iaddr),
    .io_trace_0_insn(csr_io_trace_0_insn),
    .io_trace_0_exception(csr_io_trace_0_exception),
    .io_customCSRs_0_value(csr_io_customCSRs_0_value)
  );
  BreakpointUnit bpu (
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st)
  );
  ALU alu (
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div (
    .clock(div_clock),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  PlusArgTimeout PlusArgTimeout (
    .clock(PlusArgTimeout_clock),
    .reset(PlusArgTimeout_reset),
    .io_count(PlusArgTimeout_io_count)
  );
  assign rf_id_rs_MPORT_en = 1'h1;
  assign rf_id_rs_MPORT_addr = ~id_raddr1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rf_id_rs_MPORT_data = rf[rf_id_rs_MPORT_addr];
  `else
  assign rf_id_rs_MPORT_data = rf_id_rs_MPORT_addr >= 5'h1f ? _RAND_1[31:0] : rf[rf_id_rs_MPORT_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rf_id_rs_MPORT_1_en = 1'h1;
  assign rf_id_rs_MPORT_1_addr = ~id_raddr2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rf_id_rs_MPORT_1_data = rf[rf_id_rs_MPORT_1_addr];
  `else
  assign rf_id_rs_MPORT_1_data = rf_id_rs_MPORT_1_addr >= 5'h1f ? _RAND_2[31:0] : rf[rf_id_rs_MPORT_1_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rf_MPORT_data = _rf_wdata_T ? io_dmem_resp_bits_data : _rf_wdata_T_5;
  assign rf_MPORT_addr = ~rf_waddr;
  assign rf_MPORT_mask = 1'h1;
  assign rf_MPORT_en = rf_wen & _T_139;
  assign io_imem_might_request = imem_might_request_reg;
  assign io_imem_req_valid = take_pc_wb | take_pc_mem;
  assign io_imem_req_bits_pc = wb_xcpt | csr_io_eret ? csr_io_evec : _io_imem_req_bits_pc_T_1;
  assign io_imem_req_bits_speculative = ~take_pc_wb;
  assign io_imem_sfence_valid = wb_reg_valid & wb_reg_sfence;
  assign io_imem_sfence_bits_rs1 = wb_reg_mem_size[0];
  assign io_imem_sfence_bits_rs2 = wb_reg_mem_size[1];
  assign io_imem_sfence_bits_addr = wb_reg_wdata;
  assign io_imem_resp_ready = ibuf_io_imem_ready;
  assign io_imem_btb_update_valid = mem_reg_valid & _wb_reg_replay_T & mem_wrong_npc & (~mem_cfi | mem_cfi_taken);
  assign io_imem_btb_update_bits_prediction_entry = mem_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_pc = ~_io_imem_btb_update_bits_pc_T_1;
  assign io_imem_btb_update_bits_isValid = mem_ctrl_branch | mem_ctrl_jalr | mem_ctrl_jal;
  assign io_imem_btb_update_bits_br_pc = mem_reg_pc + _GEN_256;
  assign io_imem_btb_update_bits_cfiType = (mem_ctrl_jal | mem_ctrl_jalr) & mem_waddr[0] ? 2'h2 :
    _io_imem_btb_update_bits_cfiType_T_10;
  assign io_imem_bht_update_valid = mem_reg_valid & _wb_reg_replay_T;
  assign io_imem_bht_update_bits_prediction_history = mem_reg_btb_resp_bht_history;
  assign io_imem_bht_update_bits_pc = io_imem_btb_update_bits_pc;
  assign io_imem_bht_update_bits_branch = mem_ctrl_branch;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_mispredict = ex_pc_valid ? mem_npc != ex_reg_pc : _mem_wrong_npc_T_3;
  assign io_imem_flush_icache = wb_reg_valid & wb_ctrl_fence_i & ~io_dmem_s2_nack;
  assign io_imem_progress = io_imem_progress_REG;
  assign io_dmem_req_valid = ex_reg_valid & ex_ctrl_mem;
  assign io_dmem_req_bits_addr = alu_io_adder_out;
  assign io_dmem_req_bits_tag = {{1'd0}, ex_dcache_tag};
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_size = ex_reg_mem_size;
  assign io_dmem_req_bits_signed = ~ex_reg_inst[14];
  assign io_dmem_req_bits_dprv = csr_io_status_dprv;
  assign io_dmem_req_bits_dv = 1'h0;
  assign io_dmem_s1_kill = killm_common | mem_ldst_xcpt | fpu_kill_mem;
  assign io_dmem_s1_data_data = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign io_ptw_ptbr_mode = csr_io_ptbr_mode;
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn;
  assign io_ptw_sfence_valid = io_imem_sfence_valid;
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1;
  assign io_ptw_status_debug = csr_io_status_debug;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_mxr = csr_io_status_mxr;
  assign io_ptw_status_sum = csr_io_status_sum;
  assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l;
  assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a;
  assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x;
  assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w;
  assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r;
  assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr;
  assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask;
  assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l;
  assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a;
  assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x;
  assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w;
  assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r;
  assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr;
  assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask;
  assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l;
  assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a;
  assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x;
  assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w;
  assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r;
  assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr;
  assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask;
  assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l;
  assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a;
  assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x;
  assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w;
  assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r;
  assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr;
  assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask;
  assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l;
  assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a;
  assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x;
  assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w;
  assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r;
  assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr;
  assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask;
  assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l;
  assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a;
  assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x;
  assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w;
  assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r;
  assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr;
  assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask;
  assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l;
  assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a;
  assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x;
  assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w;
  assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r;
  assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr;
  assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask;
  assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l;
  assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a;
  assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x;
  assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w;
  assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r;
  assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr;
  assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask;
  assign io_ptw_customCSRs_csrs_0_value = csr_io_customCSRs_0_value;
  assign io_fpu_inst = ibuf_io_inst_0_bits_inst_bits;
  assign io_fpu_fromint_data = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6;
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_dmem_resp_val = dmem_resp_valid & io_dmem_resp_bits_tag[0];
  assign io_fpu_dmem_resp_tag = io_dmem_resp_bits_tag[5:1];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_valid = _ex_reg_valid_T & id_ctrl_decoder_1;
  assign io_fpu_killx = take_pc_mem_wb | replay_ex | ~ex_reg_valid;
  assign io_fpu_killm = dcache_kill_mem | take_pc_wb | mem_reg_xcpt | ~mem_reg_valid;
  assign io_rocc_cmd_valid = replay_wb_rocc & _io_imem_progress_T;
  assign io_wfi = csr_io_status_wfi;
  assign ibuf_clock = clock;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid;
  assign ibuf_io_imem_bits_btb_taken = io_imem_resp_bits_btb_taken;
  assign ibuf_io_imem_bits_btb_bridx = io_imem_resp_bits_btb_bridx;
  assign ibuf_io_imem_bits_btb_entry = io_imem_resp_bits_btb_entry;
  assign ibuf_io_imem_bits_btb_bht_history = io_imem_resp_bits_btb_bht_history;
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc;
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data;
  assign ibuf_io_imem_bits_xcpt_pf_inst = io_imem_resp_bits_xcpt_pf_inst;
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst;
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay;
  assign ibuf_io_kill = take_pc_wb | take_pc_mem;
  assign ibuf_io_inst_0_ready = ~ctrl_stalld;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_ungated_clock = clock;
  assign csr_io_interrupts_debug = io_interrupts_debug;
  assign csr_io_interrupts_mtip = io_interrupts_mtip;
  assign csr_io_interrupts_msip = io_interrupts_msip;
  assign csr_io_interrupts_meip = io_interrupts_meip;
  assign csr_io_interrupts_seip = io_interrupts_seip;
  assign csr_io_hartid = io_hartid;
  assign csr_io_rw_addr = wb_reg_inst[31:20];
  assign csr_io_rw_cmd = wb_ctrl_csr & _csr_io_rw_cmd_T_1;
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_decode_0_inst = ibuf_io_inst_0_bits_inst_bits;
  assign csr_io_exception = wb_reg_xcpt | _T_97 | _T_99 | _T_105 | _T_107 | _T_109 | _T_111;
  assign csr_io_retire = wb_reg_valid & ~replay_wb & ~wb_xcpt;
  assign csr_io_cause = wb_reg_xcpt ? wb_reg_cause : {{27'd0}, _T_125};
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_tval = tval_valid ? wb_reg_wdata : 32'h0;
  assign csr_io_gva = wb_xcpt & (tval_dmem_addr & wb_reg_hls_or_dv);
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid;
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits;
  assign csr_io_inst_0 = {_csr_io_inst_0_T_3,wb_reg_raw_inst[15:0]};
  assign bpu_io_status_debug = csr_io_status_debug;
  assign bpu_io_status_prv = csr_io_status_prv;
  assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action;
  assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch;
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m;
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s;
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u;
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
  assign bpu_io_bp_0_address = csr_io_bp_0_address;
  assign bpu_io_pc = ibuf_io_pc;
  assign bpu_io_ea = mem_reg_wdata;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign alu_io_in2 = 2'h1 == ex_ctrl_sel_alu2 ? $signed({{28{_ex_op2_T_1[3]}},_ex_op2_T_1}) : $signed(_ex_op2_T_5);
  assign alu_io_in1 = 2'h2 == ex_ctrl_sel_alu1 ? $signed(ex_reg_pc) : $signed(_ex_op1_T_3);
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_req_valid = ex_reg_valid & ex_ctrl_div;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_in1 = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6;
  assign div_io_req_bits_in2 = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13;
  assign div_io_req_bits_tag = ex_reg_inst[11:7];
  assign div_io_kill = killm_common & div_io_kill_REG;
  assign div_io_resp_ready = dmem_resp_replay & dmem_resp_xpu ? 1'h0 : _ctrl_stalld_T_17;
  assign PlusArgTimeout_clock = clock;
  assign PlusArgTimeout_reset = reset;
  assign PlusArgTimeout_io_count = csr_io_time;
  always @(posedge clock) begin
    if (rf_MPORT_en & rf_MPORT_mask) begin
      rf[rf_MPORT_addr] <= rf_MPORT_data;
    end
    if (unpause) begin
      id_reg_pause <= 1'h0;
    end else if (_ex_reg_valid_T) begin
      id_reg_pause <= _GEN_1;
    end
    imem_might_request_reg <= ex_pc_valid | mem_pc_valid | io_ptw_customCSRs_csrs_0_value[1];
    if (_ex_reg_valid_T) begin
      ex_ctrl_fp <= id_ctrl_decoder_1;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_rocc <= id_ctrl_decoder_2;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_branch <= id_ctrl_decoder_3;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_jal <= id_ctrl_decoder_4;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_jalr <= id_ctrl_decoder_5;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_rxs2 <= id_ctrl_decoder_6;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_rxs1 <= id_ctrl_decoder_7;
    end
    if (_ex_reg_valid_T) begin
      if (id_xcpt) begin
        if (bpu_io_xcpt_if | _T_39) begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end else if (|_T_37) begin
          ex_ctrl_sel_alu2 <= 2'h1;
        end else begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end
      end else begin
        ex_ctrl_sel_alu2 <= id_ctrl_decoder_9;
      end
    end
    if (_ex_reg_valid_T) begin
      if (id_xcpt) begin
        if (bpu_io_xcpt_if | _T_39) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else if (|_T_37) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else begin
          ex_ctrl_sel_alu1 <= 2'h1;
        end
      end else begin
        ex_ctrl_sel_alu1 <= id_ctrl_decoder_10;
      end
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_sel_imm <= id_ctrl_decoder_11;
    end
    if (_ex_reg_valid_T) begin
      if (id_xcpt) begin
        ex_ctrl_alu_fn <= 4'h0;
      end else begin
        ex_ctrl_alu_fn <= id_ctrl_decoder_13;
      end
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_mem <= id_ctrl_decoder_14;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_mem_cmd <= id_ctrl_decoder_15;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_rfs1 <= id_ctrl_decoder_16;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_rfs2 <= id_ctrl_decoder_17;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_wfd <= id_ctrl_decoder_19;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_mul <= id_ctrl_decoder_20;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_div <= id_ctrl_decoder_21;
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_wxd <= id_ctrl_decoder_22;
    end
    if (_ex_reg_valid_T) begin
      if (id_system_insn & id_ctrl_decoder_14) begin
        ex_ctrl_csr <= 3'h0;
      end else if (id_csr_ren) begin
        ex_ctrl_csr <= 3'h2;
      end else begin
        ex_ctrl_csr <= id_ctrl_decoder_23;
      end
    end
    if (_ex_reg_valid_T) begin
      ex_ctrl_fence_i <= id_ctrl_decoder_24;
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rocc <= ex_ctrl_rocc;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rxs2 <= ex_ctrl_rxs2;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rxs1 <= ex_ctrl_rxs1;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rfs1 <= ex_ctrl_rfs1;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_rfs2 <= ex_ctrl_rfs2;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_mul <= ex_ctrl_mul;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fence_i <= _GEN_80;
      end
    end
    if (mem_pc_valid) begin
      wb_ctrl_rocc <= mem_ctrl_rocc;
    end
    if (mem_pc_valid) begin
      wb_ctrl_rxs2 <= mem_ctrl_rxs2;
    end
    if (mem_pc_valid) begin
      wb_ctrl_rxs1 <= mem_ctrl_rxs1;
    end
    if (mem_pc_valid) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if (mem_pc_valid) begin
      wb_ctrl_rfs1 <= mem_ctrl_rfs1;
    end
    if (mem_pc_valid) begin
      wb_ctrl_rfs2 <= mem_ctrl_rfs2;
    end
    if (mem_pc_valid) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if (mem_pc_valid) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if (mem_pc_valid) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if (mem_pc_valid) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if (mem_pc_valid) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    ex_reg_xcpt_interrupt <= _ex_reg_replay_T_1 & csr_io_interrupt;
    ex_reg_valid <= ~ctrl_killd;
    if (_ex_reg_valid_T) begin
      if (id_xcpt) begin
        ex_reg_rvc <= _GEN_5;
      end else begin
        ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
      end
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin
      ex_reg_btb_resp_entry <= ibuf_io_btb_resp_entry;
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin
      ex_reg_btb_resp_bht_history <= ibuf_io_btb_resp_bht_history;
    end
    ex_reg_xcpt <= _ex_reg_valid_T & id_xcpt;
    if (_ex_reg_valid_T) begin
      ex_reg_flush_pipe <= id_ctrl_decoder_24 | id_csr_flush;
    end
    if (_ex_reg_valid_T) begin
      ex_reg_load_use <= id_load_use;
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin
      if (csr_io_interrupt) begin
        ex_reg_cause <= csr_io_interrupt_cause;
      end else begin
        ex_reg_cause <= {{27'd0}, _T_18};
      end
    end
    ex_reg_replay <= ~take_pc_mem_wb & ibuf_io_inst_0_valid & ibuf_io_inst_0_bits_replay;
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin
      ex_reg_pc <= ibuf_io_pc;
    end
    if (_ex_reg_valid_T) begin
      if (id_ctrl_decoder_24) begin
        ex_reg_mem_size <= 2'h0;
      end else if (_T_48) begin
        ex_reg_mem_size <= _ex_reg_mem_size_T_6;
      end else begin
        ex_reg_mem_size <= ibuf_io_inst_0_bits_inst_bits[13:12];
      end
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin
      ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin
      ex_reg_raw_inst <= ibuf_io_inst_0_bits_raw;
    end
    mem_reg_xcpt_interrupt <= _ex_reg_replay_T & ex_reg_xcpt_interrupt;
    mem_reg_valid <= ~ctrl_killx;
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_rvc <= ex_reg_rvc;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
      end
    end
    mem_reg_xcpt <= _mem_reg_valid_T & ex_xcpt;
    mem_reg_replay <= _ex_reg_replay_T & replay_ex;
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_flush_pipe <= _GEN_81;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_cause <= ex_reg_cause;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_load <= ex_ctrl_mem & _mem_reg_load_T_24;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_store <= ex_ctrl_mem & _mem_reg_store_T_22;
      end
    end
    if (mem_reg_valid & mem_reg_flush_pipe) begin
      mem_reg_sfence <= 1'h0;
    end else if (ex_pc_valid) begin
      mem_reg_sfence <= ex_sfence;
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_mem_size <= ex_reg_mem_size;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_hls_or_dv <= io_dmem_req_bits_dv;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_raw_inst <= ex_reg_raw_inst;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_reg_wdata <= _mem_reg_wdata_T;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        if (ex_ctrl_rxs2 & (ex_ctrl_mem | ex_ctrl_rocc | ex_sfence)) begin
          if (size == 2'h0) begin
            mem_reg_rs2 <= _mem_reg_rs2_T_3;
          end else begin
            mem_reg_rs2 <= _mem_reg_rs2_T_7;
          end
        end
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin
      if (ex_pc_valid) begin
        mem_br_taken <= alu_io_cmp_out;
      end
    end
    wb_reg_valid <= ~ctrl_killm;
    wb_reg_xcpt <= mem_xcpt & _wb_reg_replay_T;
    wb_reg_replay <= replay_mem & ~take_pc_wb;
    wb_reg_flush_pipe <= _wb_reg_valid_T & mem_reg_flush_pipe;
    if (mem_pc_valid) begin
      if (_T_74) begin
        wb_reg_cause <= mem_reg_cause;
      end else begin
        wb_reg_cause <= {{28'd0}, _T_78};
      end
    end
    if (mem_pc_valid) begin
      wb_reg_sfence <= mem_reg_sfence;
    end
    if (mem_pc_valid) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if (mem_pc_valid) begin
      wb_reg_mem_size <= mem_reg_mem_size;
    end
    if (mem_pc_valid) begin
      wb_reg_hls_or_dv <= mem_reg_hls_or_dv;
    end
    if (mem_pc_valid) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if (mem_pc_valid) begin
      wb_reg_raw_inst <= mem_reg_raw_inst;
    end
    if (mem_pc_valid) begin
      if (_take_pc_mem_T & mem_ctrl_fp & mem_ctrl_wxd) begin
        wb_reg_wdata <= io_fpu_toint_data;
      end else begin
        wb_reg_wdata <= mem_int_wdata;
      end
    end
    if (reset) begin
      id_reg_fence <= 1'h0;
    end else if (_ex_reg_valid_T) begin
      id_reg_fence <= _GEN_2;
    end else if (~id_mem_busy) begin
      id_reg_fence <= 1'h0;
    end
    if (_ex_reg_valid_T) begin
      if (id_illegal_insn) begin
        ex_reg_rs_bypass_0 <= 1'h0;
      end else begin
        ex_reg_rs_bypass_0 <= do_bypass;
      end
    end
    if (_ex_reg_valid_T) begin
      ex_reg_rs_bypass_1 <= do_bypass_1;
    end
    if (_ex_reg_valid_T) begin
      if (id_illegal_insn) begin
        ex_reg_rs_lsb_0 <= inst[1:0];
      end else if (id_ctrl_decoder_7 & ~do_bypass) begin
        ex_reg_rs_lsb_0 <= id_rs_0[1:0];
      end else if (id_bypass_src_0_0) begin
        ex_reg_rs_lsb_0 <= 2'h0;
      end else begin
        ex_reg_rs_lsb_0 <= _bypass_src_T_1;
      end
    end
    if (_ex_reg_valid_T) begin
      if (id_ctrl_decoder_6 & ~do_bypass_1) begin
        ex_reg_rs_lsb_1 <= id_rs_1[1:0];
      end else if (id_bypass_src_1_0) begin
        ex_reg_rs_lsb_1 <= 2'h0;
      end else if (id_bypass_src_1_1) begin
        ex_reg_rs_lsb_1 <= 2'h1;
      end else begin
        ex_reg_rs_lsb_1 <= _bypass_src_T_2;
      end
    end
    if (_ex_reg_valid_T) begin
      if (id_illegal_insn) begin
        ex_reg_rs_msb_0 <= inst[31:2];
      end else if (id_ctrl_decoder_7 & ~do_bypass) begin
        ex_reg_rs_msb_0 <= id_rs_0[31:2];
      end
    end
    if (_ex_reg_valid_T) begin
      if (id_ctrl_decoder_6 & ~do_bypass_1) begin
        ex_reg_rs_msb_1 <= id_rs_1[31:2];
      end
    end
    if (reset) begin
      _r <= 32'h0;
    end else if (_T_159) begin
      _r <= _T_158;
    end else if (ll_wen) begin
      _r <= _T_153;
    end
    if (reset) begin
      id_stall_fpu__r <= 32'h0;
    end else if (_id_stall_fpu_T_17) begin
      id_stall_fpu__r <= _id_stall_fpu_T_16;
    end else if (_id_stall_fpu_T_12) begin
      id_stall_fpu__r <= _id_stall_fpu_T_11;
    end else if (_id_stall_fpu_T_2) begin
      id_stall_fpu__r <= _id_stall_fpu_T_5;
    end
    blocked <= _replay_ex_structural_T & _dcache_blocked_T & (blocked | io_dmem_req_valid | io_dmem_s2_nack);
    rocc_blocked <= _wb_valid_T_2 & (io_rocc_cmd_valid | rocc_blocked);
    div_io_kill_REG <= div_io_req_ready & div_io_req_valid;
    io_imem_progress_REG <= wb_reg_valid & ~replay_wb_common;
    if (ex_reg_rs_bypass_0) begin
      if (ex_reg_rs_lsb_0 == 2'h3) begin
        coreMonitorBundle_rd0val_x23 <= io_dmem_resp_bits_data_word_bypass;
      end else if (ex_reg_rs_lsb_0 == 2'h2) begin
        coreMonitorBundle_rd0val_x23 <= wb_reg_wdata;
      end else if (ex_reg_rs_lsb_0 == 2'h1) begin
        coreMonitorBundle_rd0val_x23 <= mem_reg_wdata;
      end else begin
        coreMonitorBundle_rd0val_x23 <= 32'h0;
      end
    end else begin
      coreMonitorBundle_rd0val_x23 <= _ex_rs_T_6;
    end
    coreMonitorBundle_rd0val_REG <= coreMonitorBundle_rd0val_x23;
    if (ex_reg_rs_bypass_1) begin
      if (ex_reg_rs_lsb_1 == 2'h3) begin
        coreMonitorBundle_rd1val_x29 <= io_dmem_resp_bits_data_word_bypass;
      end else if (ex_reg_rs_lsb_1 == 2'h2) begin
        coreMonitorBundle_rd1val_x29 <= wb_reg_wdata;
      end else if (ex_reg_rs_lsb_1 == 2'h1) begin
        coreMonitorBundle_rd1val_x29 <= mem_reg_wdata;
      end else begin
        coreMonitorBundle_rd1val_x29 <= 32'h0;
      end
    end else begin
      coreMonitorBundle_rd1val_x29 <= _ex_rs_T_13;
    end
    coreMonitorBundle_rd1val_REG <= coreMonitorBundle_rd1val_x29;
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~htval_valid_imem) & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~htval_valid_imem)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at RocketCore.scala:735 assert(!htval_valid_imem || io.imem.gpa.valid)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (csr_io_trace_0_valid & _csr_io_htval_T_3) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%x] W[r%d=%x][%d] R[r%d=%x] R[r%d=%x] inst=[%x] DASM(%x)\n",io_hartid,
            _io_fpu_time_T,coreMonitorBundle_valid,coreMonitorBundle_pc,_T_161,_T_162,coreMonitorBundle_wrenx,_T_164,
            _T_166,_T_168,_T_170,coreMonitorBundle_inst,coreMonitorBundle_inst);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    rf[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  id_reg_pause = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  imem_might_request_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ex_ctrl_fp = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ex_ctrl_rocc = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ex_ctrl_branch = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ex_ctrl_jal = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ex_ctrl_jalr = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ex_ctrl_rxs2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ex_ctrl_rxs1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ex_ctrl_sel_alu2 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  ex_ctrl_sel_alu1 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  ex_ctrl_sel_imm = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  ex_ctrl_alu_fn = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  ex_ctrl_mem = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ex_ctrl_mem_cmd = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  ex_ctrl_rfs1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ex_ctrl_rfs2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ex_ctrl_wfd = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ex_ctrl_mul = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ex_ctrl_div = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ex_ctrl_wxd = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  ex_ctrl_csr = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  ex_ctrl_fence_i = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_fp = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_rocc = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_branch = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_jal = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  mem_ctrl_jalr = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  mem_ctrl_rxs2 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  mem_ctrl_rxs1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  mem_ctrl_mem = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  mem_ctrl_rfs1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  mem_ctrl_rfs2 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  mem_ctrl_wfd = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  mem_ctrl_mul = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  mem_ctrl_wxd = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  mem_ctrl_csr = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  mem_ctrl_fence_i = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  wb_ctrl_rocc = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  wb_ctrl_rxs2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  wb_ctrl_rxs1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  wb_ctrl_mem = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  wb_ctrl_rfs1 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  wb_ctrl_rfs2 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  wb_ctrl_wfd = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  wb_ctrl_div = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  wb_ctrl_wxd = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  wb_ctrl_csr = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  wb_ctrl_fence_i = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ex_reg_xcpt_interrupt = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ex_reg_valid = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ex_reg_rvc = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ex_reg_btb_resp_entry = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  ex_reg_btb_resp_bht_history = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  ex_reg_xcpt = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  ex_reg_flush_pipe = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  ex_reg_load_use = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  ex_reg_cause = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  ex_reg_replay = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  ex_reg_pc = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  ex_reg_mem_size = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  ex_reg_inst = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  ex_reg_raw_inst = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mem_reg_xcpt_interrupt = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  mem_reg_valid = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  mem_reg_rvc = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  mem_reg_btb_resp_entry = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  mem_reg_btb_resp_bht_history = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  mem_reg_xcpt = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  mem_reg_replay = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  mem_reg_flush_pipe = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  mem_reg_cause = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mem_reg_slow_bypass = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  mem_reg_load = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  mem_reg_store = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  mem_reg_sfence = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  mem_reg_pc = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mem_reg_inst = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mem_reg_mem_size = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  mem_reg_hls_or_dv = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  mem_reg_raw_inst = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mem_reg_wdata = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mem_reg_rs2 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mem_br_taken = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  wb_reg_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  wb_reg_xcpt = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  wb_reg_replay = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  wb_reg_flush_pipe = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  wb_reg_cause = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  wb_reg_sfence = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  wb_reg_pc = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  wb_reg_mem_size = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  wb_reg_hls_or_dv = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  wb_reg_inst = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  wb_reg_raw_inst = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  wb_reg_wdata = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  id_reg_fence = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  ex_reg_rs_bypass_0 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  ex_reg_rs_bypass_1 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  ex_reg_rs_lsb_0 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  ex_reg_rs_lsb_1 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  ex_reg_rs_msb_0 = _RAND_105[29:0];
  _RAND_106 = {1{`RANDOM}};
  ex_reg_rs_msb_1 = _RAND_106[29:0];
  _RAND_107 = {1{`RANDOM}};
  _r = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  id_stall_fpu__r = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  blocked = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  rocc_blocked = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  div_io_kill_REG = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  io_imem_progress_REG = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  coreMonitorBundle_rd0val_x23 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  coreMonitorBundle_rd0val_REG = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  coreMonitorBundle_rd1val_x29 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  coreMonitorBundle_rd1val_REG = _RAND_116[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule