// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_210
`define RVX_GDEF_210

`define RVX_GDEF_152 6
`define RVX_GDEF_093 8
`define RVX_GDEF_427 3
`define RVX_GDEF_335 1

`define RVX_GDEF_373 (32'h 0)
`define RVX_GDEF_075 (32'h 8)
`define RVX_GDEF_395 (32'h 10)
`define RVX_GDEF_425 (32'h 18)
`define RVX_GDEF_385 (32'h 20)
`define RVX_GDEF_000 (32'h 28)
`define RVX_GDEF_344 (32'h 30)
`define RVX_GDEF_430 (32'h 38)

`define RVX_GDEF_406 (`RVX_GDEF_373)
`define RVX_GDEF_277 (`RVX_GDEF_075)
`define RVX_GDEF_399 (`RVX_GDEF_395)
`define RVX_GDEF_162 (`RVX_GDEF_425)
`define RVX_GDEF_279 (`RVX_GDEF_385)
`define RVX_GDEF_221 (`RVX_GDEF_000)
`define RVX_GDEF_134 (`RVX_GDEF_344)
`define RVX_GDEF_434 (`RVX_GDEF_430)

`define RVX_GDEF_087 3
`define RVX_GDEF_024 0
`define RVX_GDEF_381 0
`define RVX_GDEF_160 1
`define RVX_GDEF_113 2
`define RVX_GDEF_340 3
`define RVX_GDEF_122 4
`define RVX_GDEF_022 0
`define RVX_GDEF_433 1
`define RVX_GDEF_417 2

`define RVX_GDEF_183 1
`define RVX_GDEF_273 0

`define RVX_GDEF_082 32
`define RVX_GDEF_140 0

`define RVX_GDEF_229 32
`define RVX_GDEF_401 0

`define RVX_GDEF_117 32
`define RVX_GDEF_428 0

`define RVX_GDEF_431 32
`define RVX_GDEF_050 0

`define RVX_GDEF_178 32
`define RVX_GDEF_045 0

`define RVX_GDEF_070 32
`define RVX_GDEF_179 0

`define RVX_GDEF_328 2
`define RVX_GDEF_165 0
`define RVX_GDEF_017 0
`define RVX_GDEF_329 1
`define RVX_GDEF_053 2
`define RVX_GDEF_331 3
`define RVX_GDEF_081 0
`define RVX_GDEF_415 1

`define RVX_GDEF_254 16
`define RVX_GDEF_194 0

`define RVX_GDEF_424 16
`define RVX_GDEF_069 0

`define RVX_GDEF_268 16
`define RVX_GDEF_201 0

`endif