`default_nettype wire
`include "timescale.vh"
module IntXbar(
  input   auto_int_in_0,
  input   auto_int_in_1,
  output  auto_int_out_0,
  output  auto_int_out_1
);
  assign auto_int_out_0 = auto_int_in_0;
  assign auto_int_out_1 = auto_int_in_1;
endmodule