// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_266
`define RVX_GDEF_266

`define RVX_GDEF_029 6
`define RVX_GDEF_052 8
`define RVX_GDEF_380 3
`define RVX_GDEF_392 1

`define RVX_GDEF_059 (32'h 0)
`define RVX_GDEF_291 (32'h 8)
`define RVX_GDEF_196 (32'h 10)
`define RVX_GDEF_429 (32'h 18)
`define RVX_GDEF_187 (32'h 20)

`define RVX_GDEF_274 (`RVX_GDEF_059)
`define RVX_GDEF_150 (`RVX_GDEF_291)
`define RVX_GDEF_362 (`RVX_GDEF_196)
`define RVX_GDEF_208 (`RVX_GDEF_429)
`define RVX_GDEF_146 (`RVX_GDEF_187)

`define RVX_GDEF_365 1
`define RVX_GDEF_306 0
`define RVX_GDEF_155 1
`define RVX_GDEF_186 0
`define RVX_GDEF_387 0

`define RVX_GDEF_027 32
`define RVX_GDEF_156 0

`define RVX_GDEF_095 32
`define RVX_GDEF_006 0

`define RVX_GDEF_174 32
`define RVX_GDEF_228 0

`define RVX_GDEF_151 32
`define RVX_GDEF_007 0

`define RVX_GDEF_304 32
`define RVX_GDEF_241 0

`endif