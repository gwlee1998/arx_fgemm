`default_nettype wire
`include "timescale.vh"
module TLROM(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [1:0]  auto_in_a_bits_size,
  input  [9:0]  auto_in_a_bits_source,
  input  [16:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input         auto_in_a_bits_corrupt,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [1:0]  auto_in_d_bits_size,
  output [9:0]  auto_in_d_bits_source,
  output [31:0] auto_in_d_bits_data
);
  wire  monitor_clock;
  wire  monitor_reset;
  wire  monitor_io_in_a_ready;
  wire  monitor_io_in_a_valid;
  wire [2:0] monitor_io_in_a_bits_opcode;
  wire [2:0] monitor_io_in_a_bits_param;
  wire [1:0] monitor_io_in_a_bits_size;
  wire [9:0] monitor_io_in_a_bits_source;
  wire [16:0] monitor_io_in_a_bits_address;
  wire [3:0] monitor_io_in_a_bits_mask;
  wire  monitor_io_in_a_bits_corrupt;
  wire  monitor_io_in_d_ready;
  wire  monitor_io_in_d_valid;
  wire [1:0] monitor_io_in_d_bits_size;
  wire [9:0] monitor_io_in_d_bits_source;
  wire [9:0] index = auto_in_a_bits_address[11:2];
  wire [3:0] high = auto_in_a_bits_address[15:12];
  wire [31:0] _GEN_1 = 10'h1 == index ? 32'h10041b : 32'h7c105073;
  wire [31:0] _GEN_2 = 10'h2 == index ? 32'h1f41413 : _GEN_1;
  wire [31:0] _GEN_3 = 10'h3 == index ? 32'hf1402573 : _GEN_2;
  wire [31:0] _GEN_4 = 10'h4 == index ? 32'h597 : _GEN_3;
  wire [31:0] _GEN_5 = 10'h5 == index ? 32'h7058593 : _GEN_4;
  wire [31:0] _GEN_6 = 10'h6 == index ? 32'h8402 : _GEN_5;
  wire [31:0] _GEN_7 = 10'h7 == index ? 32'h0 : _GEN_6;
  wire [31:0] _GEN_8 = 10'h8 == index ? 32'h0 : _GEN_7;
  wire [31:0] _GEN_9 = 10'h9 == index ? 32'h0 : _GEN_8;
  wire [31:0] _GEN_10 = 10'ha == index ? 32'h0 : _GEN_9;
  wire [31:0] _GEN_11 = 10'hb == index ? 32'h0 : _GEN_10;
  wire [31:0] _GEN_12 = 10'hc == index ? 32'h0 : _GEN_11;
  wire [31:0] _GEN_13 = 10'hd == index ? 32'h0 : _GEN_12;
  wire [31:0] _GEN_14 = 10'he == index ? 32'h0 : _GEN_13;
  wire [31:0] _GEN_15 = 10'hf == index ? 32'h0 : _GEN_14;
  wire [31:0] _GEN_16 = 10'h10 == index ? 32'h7c105073 : _GEN_15;
  wire [31:0] _GEN_17 = 10'h11 == index ? 32'hf1402573 : _GEN_16;
  wire [31:0] _GEN_18 = 10'h12 == index ? 32'h597 : _GEN_17;
  wire [31:0] _GEN_19 = 10'h13 == index ? 32'h3858593 : _GEN_18;
  wire [31:0] _GEN_20 = 10'h14 == index ? 32'h30405073 : _GEN_19;
  wire [31:0] _GEN_21 = 10'h15 == index ? 32'h10500073 : _GEN_20;
  wire [31:0] _GEN_22 = 10'h16 == index ? 32'hbff5 : _GEN_21;
  wire [31:0] _GEN_23 = 10'h17 == index ? 32'h0 : _GEN_22;
  wire [31:0] _GEN_24 = 10'h18 == index ? 32'h0 : _GEN_23;
  wire [31:0] _GEN_25 = 10'h19 == index ? 32'h0 : _GEN_24;
  wire [31:0] _GEN_26 = 10'h1a == index ? 32'h0 : _GEN_25;
  wire [31:0] _GEN_27 = 10'h1b == index ? 32'h0 : _GEN_26;
  wire [31:0] _GEN_28 = 10'h1c == index ? 32'h0 : _GEN_27;
  wire [31:0] _GEN_29 = 10'h1d == index ? 32'h0 : _GEN_28;
  wire [31:0] _GEN_30 = 10'h1e == index ? 32'h0 : _GEN_29;
  wire [31:0] _GEN_31 = 10'h1f == index ? 32'h0 : _GEN_30;
  wire [31:0] _GEN_32 = 10'h20 == index ? 32'hedfe0dd0 : _GEN_31;
  wire [31:0] _GEN_33 = 10'h21 == index ? 32'ha5090000 : _GEN_32;
  wire [31:0] _GEN_34 = 10'h22 == index ? 32'h38000000 : _GEN_33;
  wire [31:0] _GEN_35 = 10'h23 == index ? 32'h8c070000 : _GEN_34;
  wire [31:0] _GEN_36 = 10'h24 == index ? 32'h28000000 : _GEN_35;
  wire [31:0] _GEN_37 = 10'h25 == index ? 32'h11000000 : _GEN_36;
  wire [31:0] _GEN_38 = 10'h26 == index ? 32'h10000000 : _GEN_37;
  wire [31:0] _GEN_39 = 10'h27 == index ? 32'h0 : _GEN_38;
  wire [31:0] _GEN_40 = 10'h28 == index ? 32'h19020000 : _GEN_39;
  wire [31:0] _GEN_41 = 10'h29 == index ? 32'h54070000 : _GEN_40;
  wire [31:0] _GEN_42 = 10'h2a == index ? 32'h0 : _GEN_41;
  wire [31:0] _GEN_43 = 10'h2b == index ? 32'h0 : _GEN_42;
  wire [31:0] _GEN_44 = 10'h2c == index ? 32'h0 : _GEN_43;
  wire [31:0] _GEN_45 = 10'h2d == index ? 32'h0 : _GEN_44;
  wire [31:0] _GEN_46 = 10'h2e == index ? 32'h1000000 : _GEN_45;
  wire [31:0] _GEN_47 = 10'h2f == index ? 32'h0 : _GEN_46;
  wire [31:0] _GEN_48 = 10'h30 == index ? 32'h3000000 : _GEN_47;
  wire [31:0] _GEN_49 = 10'h31 == index ? 32'h4000000 : _GEN_48;
  wire [31:0] _GEN_50 = 10'h32 == index ? 32'h0 : _GEN_49;
  wire [31:0] _GEN_51 = 10'h33 == index ? 32'h1000000 : _GEN_50;
  wire [31:0] _GEN_52 = 10'h34 == index ? 32'h3000000 : _GEN_51;
  wire [31:0] _GEN_53 = 10'h35 == index ? 32'h4000000 : _GEN_52;
  wire [31:0] _GEN_54 = 10'h36 == index ? 32'hf000000 : _GEN_53;
  wire [31:0] _GEN_55 = 10'h37 == index ? 32'h1000000 : _GEN_54;
  wire [31:0] _GEN_56 = 10'h38 == index ? 32'h3000000 : _GEN_55;
  wire [31:0] _GEN_57 = 10'h39 == index ? 32'h21000000 : _GEN_56;
  wire [31:0] _GEN_58 = 10'h3a == index ? 32'h1b000000 : _GEN_57;
  wire [31:0] _GEN_59 = 10'h3b == index ? 32'h65657266 : _GEN_58;
  wire [31:0] _GEN_60 = 10'h3c == index ? 32'h70696863 : _GEN_59;
  wire [31:0] _GEN_61 = 10'h3d == index ? 32'h6f722c73 : _GEN_60;
  wire [31:0] _GEN_62 = 10'h3e == index ? 32'h74656b63 : _GEN_61;
  wire [31:0] _GEN_63 = 10'h3f == index ? 32'h70696863 : _GEN_62;
  wire [31:0] _GEN_64 = 10'h40 == index ? 32'h6b6e752d : _GEN_63;
  wire [31:0] _GEN_65 = 10'h41 == index ? 32'h6e776f6e : _GEN_64;
  wire [31:0] _GEN_66 = 10'h42 == index ? 32'h7665642d : _GEN_65;
  wire [31:0] _GEN_67 = 10'h43 == index ? 32'h0 : _GEN_66;
  wire [31:0] _GEN_68 = 10'h44 == index ? 32'h3000000 : _GEN_67;
  wire [31:0] _GEN_69 = 10'h45 == index ? 32'h1d000000 : _GEN_68;
  wire [31:0] _GEN_70 = 10'h46 == index ? 32'h26000000 : _GEN_69;
  wire [31:0] _GEN_71 = 10'h47 == index ? 32'h65657266 : _GEN_70;
  wire [31:0] _GEN_72 = 10'h48 == index ? 32'h70696863 : _GEN_71;
  wire [31:0] _GEN_73 = 10'h49 == index ? 32'h6f722c73 : _GEN_72;
  wire [31:0] _GEN_74 = 10'h4a == index ? 32'h74656b63 : _GEN_73;
  wire [31:0] _GEN_75 = 10'h4b == index ? 32'h70696863 : _GEN_74;
  wire [31:0] _GEN_76 = 10'h4c == index ? 32'h6b6e752d : _GEN_75;
  wire [31:0] _GEN_77 = 10'h4d == index ? 32'h6e776f6e : _GEN_76;
  wire [31:0] _GEN_78 = 10'h4e == index ? 32'h0 : _GEN_77;
  wire [31:0] _GEN_79 = 10'h4f == index ? 32'h1000000 : _GEN_78;
  wire [31:0] _GEN_80 = 10'h50 == index ? 32'h73757063 : _GEN_79;
  wire [31:0] _GEN_81 = 10'h51 == index ? 32'h0 : _GEN_80;
  wire [31:0] _GEN_82 = 10'h52 == index ? 32'h3000000 : _GEN_81;
  wire [31:0] _GEN_83 = 10'h53 == index ? 32'h4000000 : _GEN_82;
  wire [31:0] _GEN_84 = 10'h54 == index ? 32'h0 : _GEN_83;
  wire [31:0] _GEN_85 = 10'h55 == index ? 32'h1000000 : _GEN_84;
  wire [31:0] _GEN_86 = 10'h56 == index ? 32'h3000000 : _GEN_85;
  wire [31:0] _GEN_87 = 10'h57 == index ? 32'h4000000 : _GEN_86;
  wire [31:0] _GEN_88 = 10'h58 == index ? 32'hf000000 : _GEN_87;
  wire [31:0] _GEN_89 = 10'h59 == index ? 32'h0 : _GEN_88;
  wire [31:0] _GEN_90 = 10'h5a == index ? 32'h3000000 : _GEN_89;
  wire [31:0] _GEN_91 = 10'h5b == index ? 32'h4000000 : _GEN_90;
  wire [31:0] _GEN_92 = 10'h5c == index ? 32'h2c000000 : _GEN_91;
  wire [31:0] _GEN_93 = 10'h5d == index ? 32'h40420f00 : _GEN_92;
  wire [31:0] _GEN_94 = 10'h5e == index ? 32'h1000000 : _GEN_93;
  wire [31:0] _GEN_95 = 10'h5f == index ? 32'h40757063 : _GEN_94;
  wire [31:0] _GEN_96 = 10'h60 == index ? 32'h30 : _GEN_95;
  wire [31:0] _GEN_97 = 10'h61 == index ? 32'h3000000 : _GEN_96;
  wire [31:0] _GEN_98 = 10'h62 == index ? 32'h4000000 : _GEN_97;
  wire [31:0] _GEN_99 = 10'h63 == index ? 32'h3f000000 : _GEN_98;
  wire [31:0] _GEN_100 = 10'h64 == index ? 32'h0 : _GEN_99;
  wire [31:0] _GEN_101 = 10'h65 == index ? 32'h3000000 : _GEN_100;
  wire [31:0] _GEN_102 = 10'h66 == index ? 32'h15000000 : _GEN_101;
  wire [31:0] _GEN_103 = 10'h67 == index ? 32'h1b000000 : _GEN_102;
  wire [31:0] _GEN_104 = 10'h68 == index ? 32'h69666973 : _GEN_103;
  wire [31:0] _GEN_105 = 10'h69 == index ? 32'h722c6576 : _GEN_104;
  wire [31:0] _GEN_106 = 10'h6a == index ? 32'h656b636f : _GEN_105;
  wire [31:0] _GEN_107 = 10'h6b == index ? 32'h72003074 : _GEN_106;
  wire [31:0] _GEN_108 = 10'h6c == index ? 32'h76637369 : _GEN_107;
  wire [31:0] _GEN_109 = 10'h6d == index ? 32'h0 : _GEN_108;
  wire [31:0] _GEN_110 = 10'h6e == index ? 32'h3000000 : _GEN_109;
  wire [31:0] _GEN_111 = 10'h6f == index ? 32'h4000000 : _GEN_110;
  wire [31:0] _GEN_112 = 10'h70 == index ? 32'h4f000000 : _GEN_111;
  wire [31:0] _GEN_113 = 10'h71 == index ? 32'h40000000 : _GEN_112;
  wire [31:0] _GEN_114 = 10'h72 == index ? 32'h3000000 : _GEN_113;
  wire [31:0] _GEN_115 = 10'h73 == index ? 32'h4000000 : _GEN_114;
  wire [31:0] _GEN_116 = 10'h74 == index ? 32'h62000000 : _GEN_115;
  wire [31:0] _GEN_117 = 10'h75 == index ? 32'h40000000 : _GEN_116;
  wire [31:0] _GEN_118 = 10'h76 == index ? 32'h3000000 : _GEN_117;
  wire [31:0] _GEN_119 = 10'h77 == index ? 32'h4000000 : _GEN_118;
  wire [31:0] _GEN_120 = 10'h78 == index ? 32'h6f000000 : _GEN_119;
  wire [31:0] _GEN_121 = 10'h79 == index ? 32'h400000 : _GEN_120;
  wire [31:0] _GEN_122 = 10'h7a == index ? 32'h3000000 : _GEN_121;
  wire [31:0] _GEN_123 = 10'h7b == index ? 32'h4000000 : _GEN_122;
  wire [31:0] _GEN_124 = 10'h7c == index ? 32'h7c000000 : _GEN_123;
  wire [31:0] _GEN_125 = 10'h7d == index ? 32'h1000000 : _GEN_124;
  wire [31:0] _GEN_126 = 10'h7e == index ? 32'h3000000 : _GEN_125;
  wire [31:0] _GEN_127 = 10'h7f == index ? 32'h4000000 : _GEN_126;
  wire [31:0] _GEN_128 = 10'h80 == index ? 32'h87000000 : _GEN_127;
  wire [31:0] _GEN_129 = 10'h81 == index ? 32'h20000000 : _GEN_128;
  wire [31:0] _GEN_130 = 10'h82 == index ? 32'h3000000 : _GEN_129;
  wire [31:0] _GEN_131 = 10'h83 == index ? 32'h4000000 : _GEN_130;
  wire [31:0] _GEN_132 = 10'h84 == index ? 32'h92000000 : _GEN_131;
  wire [31:0] _GEN_133 = 10'h85 == index ? 32'h757063 : _GEN_132;
  wire [31:0] _GEN_134 = 10'h86 == index ? 32'h3000000 : _GEN_133;
  wire [31:0] _GEN_135 = 10'h87 == index ? 32'h4000000 : _GEN_134;
  wire [31:0] _GEN_136 = 10'h88 == index ? 32'h9e000000 : _GEN_135;
  wire [31:0] _GEN_137 = 10'h89 == index ? 32'h1000000 : _GEN_136;
  wire [31:0] _GEN_138 = 10'h8a == index ? 32'h3000000 : _GEN_137;
  wire [31:0] _GEN_139 = 10'h8b == index ? 32'h4000000 : _GEN_138;
  wire [31:0] _GEN_140 = 10'h8c == index ? 32'hbd000000 : _GEN_139;
  wire [31:0] _GEN_141 = 10'h8d == index ? 32'h40000000 : _GEN_140;
  wire [31:0] _GEN_142 = 10'h8e == index ? 32'h3000000 : _GEN_141;
  wire [31:0] _GEN_143 = 10'h8f == index ? 32'h4000000 : _GEN_142;
  wire [31:0] _GEN_144 = 10'h90 == index ? 32'hd0000000 : _GEN_143;
  wire [31:0] _GEN_145 = 10'h91 == index ? 32'h40000000 : _GEN_144;
  wire [31:0] _GEN_146 = 10'h92 == index ? 32'h3000000 : _GEN_145;
  wire [31:0] _GEN_147 = 10'h93 == index ? 32'h4000000 : _GEN_146;
  wire [31:0] _GEN_148 = 10'h94 == index ? 32'hdd000000 : _GEN_147;
  wire [31:0] _GEN_149 = 10'h95 == index ? 32'h400000 : _GEN_148;
  wire [31:0] _GEN_150 = 10'h96 == index ? 32'h3000000 : _GEN_149;
  wire [31:0] _GEN_151 = 10'h97 == index ? 32'h4000000 : _GEN_150;
  wire [31:0] _GEN_152 = 10'h98 == index ? 32'hea000000 : _GEN_151;
  wire [31:0] _GEN_153 = 10'h99 == index ? 32'h1000000 : _GEN_152;
  wire [31:0] _GEN_154 = 10'h9a == index ? 32'h3000000 : _GEN_153;
  wire [31:0] _GEN_155 = 10'h9b == index ? 32'h4000000 : _GEN_154;
  wire [31:0] _GEN_156 = 10'h9c == index ? 32'hf5000000 : _GEN_155;
  wire [31:0] _GEN_157 = 10'h9d == index ? 32'h20000000 : _GEN_156;
  wire [31:0] _GEN_158 = 10'h9e == index ? 32'h3000000 : _GEN_157;
  wire [31:0] _GEN_159 = 10'h9f == index ? 32'hb000000 : _GEN_158;
  wire [31:0] _GEN_160 = 10'ha0 == index ? 32'h10000 : _GEN_159;
  wire [31:0] _GEN_161 = 10'ha1 == index ? 32'h63736972 : _GEN_160;
  wire [31:0] _GEN_162 = 10'ha2 == index ? 32'h76732c76 : _GEN_161;
  wire [31:0] _GEN_163 = 10'ha3 == index ? 32'h3233 : _GEN_162;
  wire [31:0] _GEN_164 = 10'ha4 == index ? 32'h3000000 : _GEN_163;
  wire [31:0] _GEN_165 = 10'ha5 == index ? 32'h8000000 : _GEN_164;
  wire [31:0] _GEN_166 = 10'ha6 == index ? 32'h9010000 : _GEN_165;
  wire [31:0] _GEN_167 = 10'ha7 == index ? 32'h1000000 : _GEN_166;
  wire [31:0] _GEN_168 = 10'ha8 == index ? 32'h2000000 : _GEN_167;
  wire [31:0] _GEN_169 = 10'ha9 == index ? 32'h3000000 : _GEN_168;
  wire [31:0] _GEN_170 = 10'haa == index ? 32'h4000000 : _GEN_169;
  wire [31:0] _GEN_171 = 10'hab == index ? 32'h1a010000 : _GEN_170;
  wire [31:0] _GEN_172 = 10'hac == index ? 32'h0 : _GEN_171;
  wire [31:0] _GEN_173 = 10'had == index ? 32'h3000000 : _GEN_172;
  wire [31:0] _GEN_174 = 10'hae == index ? 32'ha000000 : _GEN_173;
  wire [31:0] _GEN_175 = 10'haf == index ? 32'h1e010000 : _GEN_174;
  wire [31:0] _GEN_176 = 10'hb0 == index ? 32'h32337672 : _GEN_175;
  wire [31:0] _GEN_177 = 10'hb1 == index ? 32'h66616d69 : _GEN_176;
  wire [31:0] _GEN_178 = 10'hb2 == index ? 32'h63 : _GEN_177;
  wire [31:0] _GEN_179 = 10'hb3 == index ? 32'h3000000 : _GEN_178;
  wire [31:0] _GEN_180 = 10'hb4 == index ? 32'h4000000 : _GEN_179;
  wire [31:0] _GEN_181 = 10'hb5 == index ? 32'h28010000 : _GEN_180;
  wire [31:0] _GEN_182 = 10'hb6 == index ? 32'h4000000 : _GEN_181;
  wire [31:0] _GEN_183 = 10'hb7 == index ? 32'h3000000 : _GEN_182;
  wire [31:0] _GEN_184 = 10'hb8 == index ? 32'h4000000 : _GEN_183;
  wire [31:0] _GEN_185 = 10'hb9 == index ? 32'h3d010000 : _GEN_184;
  wire [31:0] _GEN_186 = 10'hba == index ? 32'h8000000 : _GEN_185;
  wire [31:0] _GEN_187 = 10'hbb == index ? 32'h3000000 : _GEN_186;
  wire [31:0] _GEN_188 = 10'hbc == index ? 32'h5000000 : _GEN_187;
  wire [31:0] _GEN_189 = 10'hbd == index ? 32'h4e010000 : _GEN_188;
  wire [31:0] _GEN_190 = 10'hbe == index ? 32'h79616b6f : _GEN_189;
  wire [31:0] _GEN_191 = 10'hbf == index ? 32'h0 : _GEN_190;
  wire [31:0] _GEN_192 = 10'hc0 == index ? 32'h3000000 : _GEN_191;
  wire [31:0] _GEN_193 = 10'hc1 == index ? 32'h4000000 : _GEN_192;
  wire [31:0] _GEN_194 = 10'hc2 == index ? 32'h2c000000 : _GEN_193;
  wire [31:0] _GEN_195 = 10'hc3 == index ? 32'h40420f00 : _GEN_194;
  wire [31:0] _GEN_196 = 10'hc4 == index ? 32'h3000000 : _GEN_195;
  wire [31:0] _GEN_197 = 10'hc5 == index ? 32'h0 : _GEN_196;
  wire [31:0] _GEN_198 = 10'hc6 == index ? 32'h55010000 : _GEN_197;
  wire [31:0] _GEN_199 = 10'hc7 == index ? 32'h1000000 : _GEN_198;
  wire [31:0] _GEN_200 = 10'hc8 == index ? 32'h65746e69 : _GEN_199;
  wire [31:0] _GEN_201 = 10'hc9 == index ? 32'h70757272 : _GEN_200;
  wire [31:0] _GEN_202 = 10'hca == index ? 32'h6f632d74 : _GEN_201;
  wire [31:0] _GEN_203 = 10'hcb == index ? 32'h6f72746e : _GEN_202;
  wire [31:0] _GEN_204 = 10'hcc == index ? 32'h72656c6c : _GEN_203;
  wire [31:0] _GEN_205 = 10'hcd == index ? 32'h0 : _GEN_204;
  wire [31:0] _GEN_206 = 10'hce == index ? 32'h3000000 : _GEN_205;
  wire [31:0] _GEN_207 = 10'hcf == index ? 32'h4000000 : _GEN_206;
  wire [31:0] _GEN_208 = 10'hd0 == index ? 32'h5f010000 : _GEN_207;
  wire [31:0] _GEN_209 = 10'hd1 == index ? 32'h1000000 : _GEN_208;
  wire [31:0] _GEN_210 = 10'hd2 == index ? 32'h3000000 : _GEN_209;
  wire [31:0] _GEN_211 = 10'hd3 == index ? 32'hf000000 : _GEN_210;
  wire [31:0] _GEN_212 = 10'hd4 == index ? 32'h1b000000 : _GEN_211;
  wire [31:0] _GEN_213 = 10'hd5 == index ? 32'h63736972 : _GEN_212;
  wire [31:0] _GEN_214 = 10'hd6 == index ? 32'h70632c76 : _GEN_213;
  wire [31:0] _GEN_215 = 10'hd7 == index ? 32'h6e692d75 : _GEN_214;
  wire [31:0] _GEN_216 = 10'hd8 == index ? 32'h6374 : _GEN_215;
  wire [31:0] _GEN_217 = 10'hd9 == index ? 32'h3000000 : _GEN_216;
  wire [31:0] _GEN_218 = 10'hda == index ? 32'h0 : _GEN_217;
  wire [31:0] _GEN_219 = 10'hdb == index ? 32'h70010000 : _GEN_218;
  wire [31:0] _GEN_220 = 10'hdc == index ? 32'h3000000 : _GEN_219;
  wire [31:0] _GEN_221 = 10'hdd == index ? 32'h4000000 : _GEN_220;
  wire [31:0] _GEN_222 = 10'hde == index ? 32'h85010000 : _GEN_221;
  wire [31:0] _GEN_223 = 10'hdf == index ? 32'h3000000 : _GEN_222;
  wire [31:0] _GEN_224 = 10'he0 == index ? 32'h2000000 : _GEN_223;
  wire [31:0] _GEN_225 = 10'he1 == index ? 32'h2000000 : _GEN_224;
  wire [31:0] _GEN_226 = 10'he2 == index ? 32'h2000000 : _GEN_225;
  wire [31:0] _GEN_227 = 10'he3 == index ? 32'h1000000 : _GEN_226;
  wire [31:0] _GEN_228 = 10'he4 == index ? 32'h6f6d656d : _GEN_227;
  wire [31:0] _GEN_229 = 10'he5 == index ? 32'h31407972 : _GEN_228;
  wire [31:0] _GEN_230 = 10'he6 == index ? 32'h30303030 : _GEN_229;
  wire [31:0] _GEN_231 = 10'he7 == index ? 32'h303030 : _GEN_230;
  wire [31:0] _GEN_232 = 10'he8 == index ? 32'h3000000 : _GEN_231;
  wire [31:0] _GEN_233 = 10'he9 == index ? 32'h7000000 : _GEN_232;
  wire [31:0] _GEN_234 = 10'hea == index ? 32'h92000000 : _GEN_233;
  wire [31:0] _GEN_235 = 10'heb == index ? 32'h6f6d656d : _GEN_234;
  wire [31:0] _GEN_236 = 10'hec == index ? 32'h7972 : _GEN_235;
  wire [31:0] _GEN_237 = 10'hed == index ? 32'h3000000 : _GEN_236;
  wire [31:0] _GEN_238 = 10'hee == index ? 32'h8000000 : _GEN_237;
  wire [31:0] _GEN_239 = 10'hef == index ? 32'h1a010000 : _GEN_238;
  wire [31:0] _GEN_240 = 10'hf0 == index ? 32'h10 : _GEN_239;
  wire [31:0] _GEN_241 = 10'hf1 == index ? 32'hb0 : _GEN_240;
  wire [31:0] _GEN_242 = 10'hf2 == index ? 32'h3000000 : _GEN_241;
  wire [31:0] _GEN_243 = 10'hf3 == index ? 32'h4000000 : _GEN_242;
  wire [31:0] _GEN_244 = 10'hf4 == index ? 32'h85010000 : _GEN_243;
  wire [31:0] _GEN_245 = 10'hf5 == index ? 32'h2000000 : _GEN_244;
  wire [31:0] _GEN_246 = 10'hf6 == index ? 32'h2000000 : _GEN_245;
  wire [31:0] _GEN_247 = 10'hf7 == index ? 32'h1000000 : _GEN_246;
  wire [31:0] _GEN_248 = 10'hf8 == index ? 32'h636f73 : _GEN_247;
  wire [31:0] _GEN_249 = 10'hf9 == index ? 32'h3000000 : _GEN_248;
  wire [31:0] _GEN_250 = 10'hfa == index ? 32'h4000000 : _GEN_249;
  wire [31:0] _GEN_251 = 10'hfb == index ? 32'h0 : _GEN_250;
  wire [31:0] _GEN_252 = 10'hfc == index ? 32'h1000000 : _GEN_251;
  wire [31:0] _GEN_253 = 10'hfd == index ? 32'h3000000 : _GEN_252;
  wire [31:0] _GEN_254 = 10'hfe == index ? 32'h4000000 : _GEN_253;
  wire [31:0] _GEN_255 = 10'hff == index ? 32'hf000000 : _GEN_254;
  wire [31:0] _GEN_256 = 10'h100 == index ? 32'h1000000 : _GEN_255;
  wire [31:0] _GEN_257 = 10'h101 == index ? 32'h3000000 : _GEN_256;
  wire [31:0] _GEN_258 = 10'h102 == index ? 32'h2c000000 : _GEN_257;
  wire [31:0] _GEN_259 = 10'h103 == index ? 32'h1b000000 : _GEN_258;
  wire [31:0] _GEN_260 = 10'h104 == index ? 32'h65657266 : _GEN_259;
  wire [31:0] _GEN_261 = 10'h105 == index ? 32'h70696863 : _GEN_260;
  wire [31:0] _GEN_262 = 10'h106 == index ? 32'h6f722c73 : _GEN_261;
  wire [31:0] _GEN_263 = 10'h107 == index ? 32'h74656b63 : _GEN_262;
  wire [31:0] _GEN_264 = 10'h108 == index ? 32'h70696863 : _GEN_263;
  wire [31:0] _GEN_265 = 10'h109 == index ? 32'h6b6e752d : _GEN_264;
  wire [31:0] _GEN_266 = 10'h10a == index ? 32'h6e776f6e : _GEN_265;
  wire [31:0] _GEN_267 = 10'h10b == index ? 32'h636f732d : _GEN_266;
  wire [31:0] _GEN_268 = 10'h10c == index ? 32'h6d697300 : _GEN_267;
  wire [31:0] _GEN_269 = 10'h10d == index ? 32'h2d656c70 : _GEN_268;
  wire [31:0] _GEN_270 = 10'h10e == index ? 32'h737562 : _GEN_269;
  wire [31:0] _GEN_271 = 10'h10f == index ? 32'h3000000 : _GEN_270;
  wire [31:0] _GEN_272 = 10'h110 == index ? 32'h0 : _GEN_271;
  wire [31:0] _GEN_273 = 10'h111 == index ? 32'h8d010000 : _GEN_272;
  wire [31:0] _GEN_274 = 10'h112 == index ? 32'h1000000 : _GEN_273;
  wire [31:0] _GEN_275 = 10'h113 == index ? 32'h6e696c63 : _GEN_274;
  wire [31:0] _GEN_276 = 10'h114 == index ? 32'h30324074 : _GEN_275;
  wire [31:0] _GEN_277 = 10'h115 == index ? 32'h30303030 : _GEN_276;
  wire [31:0] _GEN_278 = 10'h116 == index ? 32'h30 : _GEN_277;
  wire [31:0] _GEN_279 = 10'h117 == index ? 32'h3000000 : _GEN_278;
  wire [31:0] _GEN_280 = 10'h118 == index ? 32'hd000000 : _GEN_279;
  wire [31:0] _GEN_281 = 10'h119 == index ? 32'h1b000000 : _GEN_280;
  wire [31:0] _GEN_282 = 10'h11a == index ? 32'h63736972 : _GEN_281;
  wire [31:0] _GEN_283 = 10'h11b == index ? 32'h6c632c76 : _GEN_282;
  wire [31:0] _GEN_284 = 10'h11c == index ? 32'h30746e69 : _GEN_283;
  wire [31:0] _GEN_285 = 10'h11d == index ? 32'h0 : _GEN_284;
  wire [31:0] _GEN_286 = 10'h11e == index ? 32'h3000000 : _GEN_285;
  wire [31:0] _GEN_287 = 10'h11f == index ? 32'h10000000 : _GEN_286;
  wire [31:0] _GEN_288 = 10'h120 == index ? 32'h94010000 : _GEN_287;
  wire [31:0] _GEN_289 = 10'h121 == index ? 32'h3000000 : _GEN_288;
  wire [31:0] _GEN_290 = 10'h122 == index ? 32'h3000000 : _GEN_289;
  wire [31:0] _GEN_291 = 10'h123 == index ? 32'h3000000 : _GEN_290;
  wire [31:0] _GEN_292 = 10'h124 == index ? 32'h7000000 : _GEN_291;
  wire [31:0] _GEN_293 = 10'h125 == index ? 32'h3000000 : _GEN_292;
  wire [31:0] _GEN_294 = 10'h126 == index ? 32'h8000000 : _GEN_293;
  wire [31:0] _GEN_295 = 10'h127 == index ? 32'h1a010000 : _GEN_294;
  wire [31:0] _GEN_296 = 10'h128 == index ? 32'h2 : _GEN_295;
  wire [31:0] _GEN_297 = 10'h129 == index ? 32'h100 : _GEN_296;
  wire [31:0] _GEN_298 = 10'h12a == index ? 32'h3000000 : _GEN_297;
  wire [31:0] _GEN_299 = 10'h12b == index ? 32'h8000000 : _GEN_298;
  wire [31:0] _GEN_300 = 10'h12c == index ? 32'ha8010000 : _GEN_299;
  wire [31:0] _GEN_301 = 10'h12d == index ? 32'h746e6f63 : _GEN_300;
  wire [31:0] _GEN_302 = 10'h12e == index ? 32'h6c6f72 : _GEN_301;
  wire [31:0] _GEN_303 = 10'h12f == index ? 32'h2000000 : _GEN_302;
  wire [31:0] _GEN_304 = 10'h130 == index ? 32'h1000000 : _GEN_303;
  wire [31:0] _GEN_305 = 10'h131 == index ? 32'h75626564 : _GEN_304;
  wire [31:0] _GEN_306 = 10'h132 == index ? 32'h6f632d67 : _GEN_305;
  wire [31:0] _GEN_307 = 10'h133 == index ? 32'h6f72746e : _GEN_306;
  wire [31:0] _GEN_308 = 10'h134 == index ? 32'h72656c6c : _GEN_307;
  wire [31:0] _GEN_309 = 10'h135 == index ? 32'h3040 : _GEN_308;
  wire [31:0] _GEN_310 = 10'h136 == index ? 32'h3000000 : _GEN_309;
  wire [31:0] _GEN_311 = 10'h137 == index ? 32'h21000000 : _GEN_310;
  wire [31:0] _GEN_312 = 10'h138 == index ? 32'h1b000000 : _GEN_311;
  wire [31:0] _GEN_313 = 10'h139 == index ? 32'h69666973 : _GEN_312;
  wire [31:0] _GEN_314 = 10'h13a == index ? 32'h642c6576 : _GEN_313;
  wire [31:0] _GEN_315 = 10'h13b == index ? 32'h67756265 : _GEN_314;
  wire [31:0] _GEN_316 = 10'h13c == index ? 32'h3331302d : _GEN_315;
  wire [31:0] _GEN_317 = 10'h13d == index ? 32'h73697200 : _GEN_316;
  wire [31:0] _GEN_318 = 10'h13e == index ? 32'h642c7663 : _GEN_317;
  wire [31:0] _GEN_319 = 10'h13f == index ? 32'h67756265 : _GEN_318;
  wire [31:0] _GEN_320 = 10'h140 == index ? 32'h3331302d : _GEN_319;
  wire [31:0] _GEN_321 = 10'h141 == index ? 32'h0 : _GEN_320;
  wire [31:0] _GEN_322 = 10'h142 == index ? 32'h3000000 : _GEN_321;
  wire [31:0] _GEN_323 = 10'h143 == index ? 32'h4000000 : _GEN_322;
  wire [31:0] _GEN_324 = 10'h144 == index ? 32'hb2010000 : _GEN_323;
  wire [31:0] _GEN_325 = 10'h145 == index ? 32'h696d64 : _GEN_324;
  wire [31:0] _GEN_326 = 10'h146 == index ? 32'h3000000 : _GEN_325;
  wire [31:0] _GEN_327 = 10'h147 == index ? 32'h8000000 : _GEN_326;
  wire [31:0] _GEN_328 = 10'h148 == index ? 32'h94010000 : _GEN_327;
  wire [31:0] _GEN_329 = 10'h149 == index ? 32'h3000000 : _GEN_328;
  wire [31:0] _GEN_330 = 10'h14a == index ? 32'hffff0000 : _GEN_329;
  wire [31:0] _GEN_331 = 10'h14b == index ? 32'h3000000 : _GEN_330;
  wire [31:0] _GEN_332 = 10'h14c == index ? 32'h8000000 : _GEN_331;
  wire [31:0] _GEN_333 = 10'h14d == index ? 32'h1a010000 : _GEN_332;
  wire [31:0] _GEN_334 = 10'h14e == index ? 32'h0 : _GEN_333;
  wire [31:0] _GEN_335 = 10'h14f == index ? 32'h100000 : _GEN_334;
  wire [31:0] _GEN_336 = 10'h150 == index ? 32'h3000000 : _GEN_335;
  wire [31:0] _GEN_337 = 10'h151 == index ? 32'h8000000 : _GEN_336;
  wire [31:0] _GEN_338 = 10'h152 == index ? 32'ha8010000 : _GEN_337;
  wire [31:0] _GEN_339 = 10'h153 == index ? 32'h746e6f63 : _GEN_338;
  wire [31:0] _GEN_340 = 10'h154 == index ? 32'h6c6f72 : _GEN_339;
  wire [31:0] _GEN_341 = 10'h155 == index ? 32'h2000000 : _GEN_340;
  wire [31:0] _GEN_342 = 10'h156 == index ? 32'h1000000 : _GEN_341;
  wire [31:0] _GEN_343 = 10'h157 == index ? 32'h6f727265 : _GEN_342;
  wire [31:0] _GEN_344 = 10'h158 == index ? 32'h65642d72 : _GEN_343;
  wire [31:0] _GEN_345 = 10'h159 == index ? 32'h65636976 : _GEN_344;
  wire [31:0] _GEN_346 = 10'h15a == index ? 32'h30303340 : _GEN_345;
  wire [31:0] _GEN_347 = 10'h15b == index ? 32'h30 : _GEN_346;
  wire [31:0] _GEN_348 = 10'h15c == index ? 32'h3000000 : _GEN_347;
  wire [31:0] _GEN_349 = 10'h15d == index ? 32'he000000 : _GEN_348;
  wire [31:0] _GEN_350 = 10'h15e == index ? 32'h1b000000 : _GEN_349;
  wire [31:0] _GEN_351 = 10'h15f == index ? 32'h69666973 : _GEN_350;
  wire [31:0] _GEN_352 = 10'h160 == index ? 32'h652c6576 : _GEN_351;
  wire [31:0] _GEN_353 = 10'h161 == index ? 32'h726f7272 : _GEN_352;
  wire [31:0] _GEN_354 = 10'h162 == index ? 32'h30 : _GEN_353;
  wire [31:0] _GEN_355 = 10'h163 == index ? 32'h3000000 : _GEN_354;
  wire [31:0] _GEN_356 = 10'h164 == index ? 32'h8000000 : _GEN_355;
  wire [31:0] _GEN_357 = 10'h165 == index ? 32'h1a010000 : _GEN_356;
  wire [31:0] _GEN_358 = 10'h166 == index ? 32'h300000 : _GEN_357;
  wire [31:0] _GEN_359 = 10'h167 == index ? 32'h100000 : _GEN_358;
  wire [31:0] _GEN_360 = 10'h168 == index ? 32'h2000000 : _GEN_359;
  wire [31:0] _GEN_361 = 10'h169 == index ? 32'h1000000 : _GEN_360;
  wire [31:0] _GEN_362 = 10'h16a == index ? 32'h65747865 : _GEN_361;
  wire [31:0] _GEN_363 = 10'h16b == index ? 32'h6c616e72 : _GEN_362;
  wire [31:0] _GEN_364 = 10'h16c == index ? 32'h746e692d : _GEN_363;
  wire [31:0] _GEN_365 = 10'h16d == index ? 32'h75727265 : _GEN_364;
  wire [31:0] _GEN_366 = 10'h16e == index ? 32'h737470 : _GEN_365;
  wire [31:0] _GEN_367 = 10'h16f == index ? 32'h3000000 : _GEN_366;
  wire [31:0] _GEN_368 = 10'h170 == index ? 32'h4000000 : _GEN_367;
  wire [31:0] _GEN_369 = 10'h171 == index ? 32'hbf010000 : _GEN_368;
  wire [31:0] _GEN_370 = 10'h172 == index ? 32'h4000000 : _GEN_369;
  wire [31:0] _GEN_371 = 10'h173 == index ? 32'h3000000 : _GEN_370;
  wire [31:0] _GEN_372 = 10'h174 == index ? 32'h8000000 : _GEN_371;
  wire [31:0] _GEN_373 = 10'h175 == index ? 32'hd0010000 : _GEN_372;
  wire [31:0] _GEN_374 = 10'h176 == index ? 32'h1000000 : _GEN_373;
  wire [31:0] _GEN_375 = 10'h177 == index ? 32'h2000000 : _GEN_374;
  wire [31:0] _GEN_376 = 10'h178 == index ? 32'h2000000 : _GEN_375;
  wire [31:0] _GEN_377 = 10'h179 == index ? 32'h1000000 : _GEN_376;
  wire [31:0] _GEN_378 = 10'h17a == index ? 32'h65746e69 : _GEN_377;
  wire [31:0] _GEN_379 = 10'h17b == index ? 32'h70757272 : _GEN_378;
  wire [31:0] _GEN_380 = 10'h17c == index ? 32'h6f632d74 : _GEN_379;
  wire [31:0] _GEN_381 = 10'h17d == index ? 32'h6f72746e : _GEN_380;
  wire [31:0] _GEN_382 = 10'h17e == index ? 32'h72656c6c : _GEN_381;
  wire [31:0] _GEN_383 = 10'h17f == index ? 32'h30306340 : _GEN_382;
  wire [31:0] _GEN_384 = 10'h180 == index ? 32'h30303030 : _GEN_383;
  wire [31:0] _GEN_385 = 10'h181 == index ? 32'h0 : _GEN_384;
  wire [31:0] _GEN_386 = 10'h182 == index ? 32'h3000000 : _GEN_385;
  wire [31:0] _GEN_387 = 10'h183 == index ? 32'h4000000 : _GEN_386;
  wire [31:0] _GEN_388 = 10'h184 == index ? 32'h5f010000 : _GEN_387;
  wire [31:0] _GEN_389 = 10'h185 == index ? 32'h1000000 : _GEN_388;
  wire [31:0] _GEN_390 = 10'h186 == index ? 32'h3000000 : _GEN_389;
  wire [31:0] _GEN_391 = 10'h187 == index ? 32'hc000000 : _GEN_390;
  wire [31:0] _GEN_392 = 10'h188 == index ? 32'h1b000000 : _GEN_391;
  wire [31:0] _GEN_393 = 10'h189 == index ? 32'h63736972 : _GEN_392;
  wire [31:0] _GEN_394 = 10'h18a == index ? 32'h6c702c76 : _GEN_393;
  wire [31:0] _GEN_395 = 10'h18b == index ? 32'h306369 : _GEN_394;
  wire [31:0] _GEN_396 = 10'h18c == index ? 32'h3000000 : _GEN_395;
  wire [31:0] _GEN_397 = 10'h18d == index ? 32'h0 : _GEN_396;
  wire [31:0] _GEN_398 = 10'h18e == index ? 32'h70010000 : _GEN_397;
  wire [31:0] _GEN_399 = 10'h18f == index ? 32'h3000000 : _GEN_398;
  wire [31:0] _GEN_400 = 10'h190 == index ? 32'h10000000 : _GEN_399;
  wire [31:0] _GEN_401 = 10'h191 == index ? 32'h94010000 : _GEN_400;
  wire [31:0] _GEN_402 = 10'h192 == index ? 32'h3000000 : _GEN_401;
  wire [31:0] _GEN_403 = 10'h193 == index ? 32'hb000000 : _GEN_402;
  wire [31:0] _GEN_404 = 10'h194 == index ? 32'h3000000 : _GEN_403;
  wire [31:0] _GEN_405 = 10'h195 == index ? 32'h9000000 : _GEN_404;
  wire [31:0] _GEN_406 = 10'h196 == index ? 32'h3000000 : _GEN_405;
  wire [31:0] _GEN_407 = 10'h197 == index ? 32'h8000000 : _GEN_406;
  wire [31:0] _GEN_408 = 10'h198 == index ? 32'h1a010000 : _GEN_407;
  wire [31:0] _GEN_409 = 10'h199 == index ? 32'hc : _GEN_408;
  wire [31:0] _GEN_410 = 10'h19a == index ? 32'h4 : _GEN_409;
  wire [31:0] _GEN_411 = 10'h19b == index ? 32'h3000000 : _GEN_410;
  wire [31:0] _GEN_412 = 10'h19c == index ? 32'h8000000 : _GEN_411;
  wire [31:0] _GEN_413 = 10'h19d == index ? 32'ha8010000 : _GEN_412;
  wire [31:0] _GEN_414 = 10'h19e == index ? 32'h746e6f63 : _GEN_413;
  wire [31:0] _GEN_415 = 10'h19f == index ? 32'h6c6f72 : _GEN_414;
  wire [31:0] _GEN_416 = 10'h1a0 == index ? 32'h3000000 : _GEN_415;
  wire [31:0] _GEN_417 = 10'h1a1 == index ? 32'h4000000 : _GEN_416;
  wire [31:0] _GEN_418 = 10'h1a2 == index ? 32'hdb010000 : _GEN_417;
  wire [31:0] _GEN_419 = 10'h1a3 == index ? 32'h3000000 : _GEN_418;
  wire [31:0] _GEN_420 = 10'h1a4 == index ? 32'h3000000 : _GEN_419;
  wire [31:0] _GEN_421 = 10'h1a5 == index ? 32'h4000000 : _GEN_420;
  wire [31:0] _GEN_422 = 10'h1a6 == index ? 32'hee010000 : _GEN_421;
  wire [31:0] _GEN_423 = 10'h1a7 == index ? 32'h2000000 : _GEN_422;
  wire [31:0] _GEN_424 = 10'h1a8 == index ? 32'h3000000 : _GEN_423;
  wire [31:0] _GEN_425 = 10'h1a9 == index ? 32'h4000000 : _GEN_424;
  wire [31:0] _GEN_426 = 10'h1aa == index ? 32'h85010000 : _GEN_425;
  wire [31:0] _GEN_427 = 10'h1ab == index ? 32'h4000000 : _GEN_426;
  wire [31:0] _GEN_428 = 10'h1ac == index ? 32'h2000000 : _GEN_427;
  wire [31:0] _GEN_429 = 10'h1ad == index ? 32'h1000000 : _GEN_428;
  wire [31:0] _GEN_430 = 10'h1ae == index ? 32'h6f696d6d : _GEN_429;
  wire [31:0] _GEN_431 = 10'h1af == index ? 32'h726f702d : _GEN_430;
  wire [31:0] _GEN_432 = 10'h1b0 == index ? 32'h78612d74 : _GEN_431;
  wire [31:0] _GEN_433 = 10'h1b1 == index ? 32'h63403469 : _GEN_432;
  wire [31:0] _GEN_434 = 10'h1b2 == index ? 32'h30303030 : _GEN_433;
  wire [31:0] _GEN_435 = 10'h1b3 == index ? 32'h303030 : _GEN_434;
  wire [31:0] _GEN_436 = 10'h1b4 == index ? 32'h3000000 : _GEN_435;
  wire [31:0] _GEN_437 = 10'h1b5 == index ? 32'h4000000 : _GEN_436;
  wire [31:0] _GEN_438 = 10'h1b6 == index ? 32'h0 : _GEN_437;
  wire [31:0] _GEN_439 = 10'h1b7 == index ? 32'h1000000 : _GEN_438;
  wire [31:0] _GEN_440 = 10'h1b8 == index ? 32'h3000000 : _GEN_439;
  wire [31:0] _GEN_441 = 10'h1b9 == index ? 32'h4000000 : _GEN_440;
  wire [31:0] _GEN_442 = 10'h1ba == index ? 32'hf000000 : _GEN_441;
  wire [31:0] _GEN_443 = 10'h1bb == index ? 32'h1000000 : _GEN_442;
  wire [31:0] _GEN_444 = 10'h1bc == index ? 32'h3000000 : _GEN_443;
  wire [31:0] _GEN_445 = 10'h1bd == index ? 32'hb000000 : _GEN_444;
  wire [31:0] _GEN_446 = 10'h1be == index ? 32'h1b000000 : _GEN_445;
  wire [31:0] _GEN_447 = 10'h1bf == index ? 32'h706d6973 : _GEN_446;
  wire [31:0] _GEN_448 = 10'h1c0 == index ? 32'h622d656c : _GEN_447;
  wire [31:0] _GEN_449 = 10'h1c1 == index ? 32'h7375 : _GEN_448;
  wire [31:0] _GEN_450 = 10'h1c2 == index ? 32'h3000000 : _GEN_449;
  wire [31:0] _GEN_451 = 10'h1c3 == index ? 32'hc000000 : _GEN_450;
  wire [31:0] _GEN_452 = 10'h1c4 == index ? 32'h8d010000 : _GEN_451;
  wire [31:0] _GEN_453 = 10'h1c5 == index ? 32'hc0 : _GEN_452;
  wire [31:0] _GEN_454 = 10'h1c6 == index ? 32'hc0 : _GEN_453;
  wire [31:0] _GEN_455 = 10'h1c7 == index ? 32'h40 : _GEN_454;
  wire [31:0] _GEN_456 = 10'h1c8 == index ? 32'h2000000 : _GEN_455;
  wire [31:0] _GEN_457 = 10'h1c9 == index ? 32'h1000000 : _GEN_456;
  wire [31:0] _GEN_458 = 10'h1ca == index ? 32'h406d6f72 : _GEN_457;
  wire [31:0] _GEN_459 = 10'h1cb == index ? 32'h30303031 : _GEN_458;
  wire [31:0] _GEN_460 = 10'h1cc == index ? 32'h30 : _GEN_459;
  wire [31:0] _GEN_461 = 10'h1cd == index ? 32'h3000000 : _GEN_460;
  wire [31:0] _GEN_462 = 10'h1ce == index ? 32'hc000000 : _GEN_461;
  wire [31:0] _GEN_463 = 10'h1cf == index ? 32'h1b000000 : _GEN_462;
  wire [31:0] _GEN_464 = 10'h1d0 == index ? 32'h69666973 : _GEN_463;
  wire [31:0] _GEN_465 = 10'h1d1 == index ? 32'h722c6576 : _GEN_464;
  wire [31:0] _GEN_466 = 10'h1d2 == index ? 32'h306d6f : _GEN_465;
  wire [31:0] _GEN_467 = 10'h1d3 == index ? 32'h3000000 : _GEN_466;
  wire [31:0] _GEN_468 = 10'h1d4 == index ? 32'h8000000 : _GEN_467;
  wire [31:0] _GEN_469 = 10'h1d5 == index ? 32'h1a010000 : _GEN_468;
  wire [31:0] _GEN_470 = 10'h1d6 == index ? 32'h100 : _GEN_469;
  wire [31:0] _GEN_471 = 10'h1d7 == index ? 32'h100 : _GEN_470;
  wire [31:0] _GEN_472 = 10'h1d8 == index ? 32'h3000000 : _GEN_471;
  wire [31:0] _GEN_473 = 10'h1d9 == index ? 32'h4000000 : _GEN_472;
  wire [31:0] _GEN_474 = 10'h1da == index ? 32'ha8010000 : _GEN_473;
  wire [31:0] _GEN_475 = 10'h1db == index ? 32'h6d656d : _GEN_474;
  wire [31:0] _GEN_476 = 10'h1dc == index ? 32'h3000000 : _GEN_475;
  wire [31:0] _GEN_477 = 10'h1dd == index ? 32'h4000000 : _GEN_476;
  wire [31:0] _GEN_478 = 10'h1de == index ? 32'h85010000 : _GEN_477;
  wire [31:0] _GEN_479 = 10'h1df == index ? 32'h1000000 : _GEN_478;
  wire [31:0] _GEN_480 = 10'h1e0 == index ? 32'h2000000 : _GEN_479;
  wire [31:0] _GEN_481 = 10'h1e1 == index ? 32'h1000000 : _GEN_480;
  wire [31:0] _GEN_482 = 10'h1e2 == index ? 32'h73627573 : _GEN_481;
  wire [31:0] _GEN_483 = 10'h1e3 == index ? 32'h65747379 : _GEN_482;
  wire [31:0] _GEN_484 = 10'h1e4 == index ? 32'h62705f6d : _GEN_483;
  wire [31:0] _GEN_485 = 10'h1e5 == index ? 32'h635f7375 : _GEN_484;
  wire [31:0] _GEN_486 = 10'h1e6 == index ? 32'h6b636f6c : _GEN_485;
  wire [31:0] _GEN_487 = 10'h1e7 == index ? 32'h0 : _GEN_486;
  wire [31:0] _GEN_488 = 10'h1e8 == index ? 32'h3000000 : _GEN_487;
  wire [31:0] _GEN_489 = 10'h1e9 == index ? 32'h4000000 : _GEN_488;
  wire [31:0] _GEN_490 = 10'h1ea == index ? 32'hf9010000 : _GEN_489;
  wire [31:0] _GEN_491 = 10'h1eb == index ? 32'h0 : _GEN_490;
  wire [31:0] _GEN_492 = 10'h1ec == index ? 32'h3000000 : _GEN_491;
  wire [31:0] _GEN_493 = 10'h1ed == index ? 32'h4000000 : _GEN_492;
  wire [31:0] _GEN_494 = 10'h1ee == index ? 32'h3f000000 : _GEN_493;
  wire [31:0] _GEN_495 = 10'h1ef == index ? 32'he1f505 : _GEN_494;
  wire [31:0] _GEN_496 = 10'h1f0 == index ? 32'h3000000 : _GEN_495;
  wire [31:0] _GEN_497 = 10'h1f1 == index ? 32'h15000000 : _GEN_496;
  wire [31:0] _GEN_498 = 10'h1f2 == index ? 32'h6020000 : _GEN_497;
  wire [31:0] _GEN_499 = 10'h1f3 == index ? 32'h73627573 : _GEN_498;
  wire [31:0] _GEN_500 = 10'h1f4 == index ? 32'h65747379 : _GEN_499;
  wire [31:0] _GEN_501 = 10'h1f5 == index ? 32'h62705f6d : _GEN_500;
  wire [31:0] _GEN_502 = 10'h1f6 == index ? 32'h635f7375 : _GEN_501;
  wire [31:0] _GEN_503 = 10'h1f7 == index ? 32'h6b636f6c : _GEN_502;
  wire [31:0] _GEN_504 = 10'h1f8 == index ? 32'h0 : _GEN_503;
  wire [31:0] _GEN_505 = 10'h1f9 == index ? 32'h3000000 : _GEN_504;
  wire [31:0] _GEN_506 = 10'h1fa == index ? 32'hc000000 : _GEN_505;
  wire [31:0] _GEN_507 = 10'h1fb == index ? 32'h1b000000 : _GEN_506;
  wire [31:0] _GEN_508 = 10'h1fc == index ? 32'h65786966 : _GEN_507;
  wire [31:0] _GEN_509 = 10'h1fd == index ? 32'h6c632d64 : _GEN_508;
  wire [31:0] _GEN_510 = 10'h1fe == index ? 32'h6b636f : _GEN_509;
  wire [31:0] _GEN_511 = 10'h1ff == index ? 32'h2000000 : _GEN_510;
  wire [31:0] _GEN_512 = 10'h200 == index ? 32'h2000000 : _GEN_511;
  wire [31:0] _GEN_513 = 10'h201 == index ? 32'h2000000 : _GEN_512;
  wire [31:0] _GEN_514 = 10'h202 == index ? 32'h9000000 : _GEN_513;
  wire [31:0] _GEN_515 = 10'h203 == index ? 32'h64646123 : _GEN_514;
  wire [31:0] _GEN_516 = 10'h204 == index ? 32'h73736572 : _GEN_515;
  wire [31:0] _GEN_517 = 10'h205 == index ? 32'h6c65632d : _GEN_516;
  wire [31:0] _GEN_518 = 10'h206 == index ? 32'h2300736c : _GEN_517;
  wire [31:0] _GEN_519 = 10'h207 == index ? 32'h657a6973 : _GEN_518;
  wire [31:0] _GEN_520 = 10'h208 == index ? 32'h6c65632d : _GEN_519;
  wire [31:0] _GEN_521 = 10'h209 == index ? 32'h6300736c : _GEN_520;
  wire [31:0] _GEN_522 = 10'h20a == index ? 32'h61706d6f : _GEN_521;
  wire [31:0] _GEN_523 = 10'h20b == index ? 32'h6c626974 : _GEN_522;
  wire [31:0] _GEN_524 = 10'h20c == index ? 32'h6f6d0065 : _GEN_523;
  wire [31:0] _GEN_525 = 10'h20d == index ? 32'h6c6564 : _GEN_524;
  wire [31:0] _GEN_526 = 10'h20e == index ? 32'h656d6974 : _GEN_525;
  wire [31:0] _GEN_527 = 10'h20f == index ? 32'h65736162 : _GEN_526;
  wire [31:0] _GEN_528 = 10'h210 == index ? 32'h6572662d : _GEN_527;
  wire [31:0] _GEN_529 = 10'h211 == index ? 32'h6e657571 : _GEN_528;
  wire [31:0] _GEN_530 = 10'h212 == index ? 32'h63007963 : _GEN_529;
  wire [31:0] _GEN_531 = 10'h213 == index ? 32'h6b636f6c : _GEN_530;
  wire [31:0] _GEN_532 = 10'h214 == index ? 32'h6572662d : _GEN_531;
  wire [31:0] _GEN_533 = 10'h215 == index ? 32'h6e657571 : _GEN_532;
  wire [31:0] _GEN_534 = 10'h216 == index ? 32'h64007963 : _GEN_533;
  wire [31:0] _GEN_535 = 10'h217 == index ? 32'h6361632d : _GEN_534;
  wire [31:0] _GEN_536 = 10'h218 == index ? 32'h622d6568 : _GEN_535;
  wire [31:0] _GEN_537 = 10'h219 == index ? 32'h6b636f6c : _GEN_536;
  wire [31:0] _GEN_538 = 10'h21a == index ? 32'h7a69732d : _GEN_537;
  wire [31:0] _GEN_539 = 10'h21b == index ? 32'h2d640065 : _GEN_538;
  wire [31:0] _GEN_540 = 10'h21c == index ? 32'h68636163 : _GEN_539;
  wire [31:0] _GEN_541 = 10'h21d == index ? 32'h65732d65 : _GEN_540;
  wire [31:0] _GEN_542 = 10'h21e == index ? 32'h64007374 : _GEN_541;
  wire [31:0] _GEN_543 = 10'h21f == index ? 32'h6361632d : _GEN_542;
  wire [31:0] _GEN_544 = 10'h220 == index ? 32'h732d6568 : _GEN_543;
  wire [31:0] _GEN_545 = 10'h221 == index ? 32'h657a69 : _GEN_544;
  wire [31:0] _GEN_546 = 10'h222 == index ? 32'h6c742d64 : _GEN_545;
  wire [31:0] _GEN_547 = 10'h223 == index ? 32'h65732d62 : _GEN_546;
  wire [31:0] _GEN_548 = 10'h224 == index ? 32'h64007374 : _GEN_547;
  wire [31:0] _GEN_549 = 10'h225 == index ? 32'h626c742d : _GEN_548;
  wire [31:0] _GEN_550 = 10'h226 == index ? 32'h7a69732d : _GEN_549;
  wire [31:0] _GEN_551 = 10'h227 == index ? 32'h65640065 : _GEN_550;
  wire [31:0] _GEN_552 = 10'h228 == index ? 32'h65636976 : _GEN_551;
  wire [31:0] _GEN_553 = 10'h229 == index ? 32'h7079745f : _GEN_552;
  wire [31:0] _GEN_554 = 10'h22a == index ? 32'h61680065 : _GEN_553;
  wire [31:0] _GEN_555 = 10'h22b == index ? 32'h61776472 : _GEN_554;
  wire [31:0] _GEN_556 = 10'h22c == index ? 32'h652d6572 : _GEN_555;
  wire [31:0] _GEN_557 = 10'h22d == index ? 32'h2d636578 : _GEN_556;
  wire [31:0] _GEN_558 = 10'h22e == index ? 32'h61657262 : _GEN_557;
  wire [31:0] _GEN_559 = 10'h22f == index ? 32'h696f706b : _GEN_558;
  wire [31:0] _GEN_560 = 10'h230 == index ? 32'h632d746e : _GEN_559;
  wire [31:0] _GEN_561 = 10'h231 == index ? 32'h746e756f : _GEN_560;
  wire [31:0] _GEN_562 = 10'h232 == index ? 32'h632d6900 : _GEN_561;
  wire [31:0] _GEN_563 = 10'h233 == index ? 32'h65686361 : _GEN_562;
  wire [31:0] _GEN_564 = 10'h234 == index ? 32'h6f6c622d : _GEN_563;
  wire [31:0] _GEN_565 = 10'h235 == index ? 32'h732d6b63 : _GEN_564;
  wire [31:0] _GEN_566 = 10'h236 == index ? 32'h657a69 : _GEN_565;
  wire [31:0] _GEN_567 = 10'h237 == index ? 32'h61632d69 : _GEN_566;
  wire [31:0] _GEN_568 = 10'h238 == index ? 32'h2d656863 : _GEN_567;
  wire [31:0] _GEN_569 = 10'h239 == index ? 32'h73746573 : _GEN_568;
  wire [31:0] _GEN_570 = 10'h23a == index ? 32'h632d6900 : _GEN_569;
  wire [31:0] _GEN_571 = 10'h23b == index ? 32'h65686361 : _GEN_570;
  wire [31:0] _GEN_572 = 10'h23c == index ? 32'h7a69732d : _GEN_571;
  wire [31:0] _GEN_573 = 10'h23d == index ? 32'h2d690065 : _GEN_572;
  wire [31:0] _GEN_574 = 10'h23e == index ? 32'h2d626c74 : _GEN_573;
  wire [31:0] _GEN_575 = 10'h23f == index ? 32'h73746573 : _GEN_574;
  wire [31:0] _GEN_576 = 10'h240 == index ? 32'h742d6900 : _GEN_575;
  wire [31:0] _GEN_577 = 10'h241 == index ? 32'h732d626c : _GEN_576;
  wire [31:0] _GEN_578 = 10'h242 == index ? 32'h657a69 : _GEN_577;
  wire [31:0] _GEN_579 = 10'h243 == index ? 32'h2d756d6d : _GEN_578;
  wire [31:0] _GEN_580 = 10'h244 == index ? 32'h65707974 : _GEN_579;
  wire [31:0] _GEN_581 = 10'h245 == index ? 32'h78656e00 : _GEN_580;
  wire [31:0] _GEN_582 = 10'h246 == index ? 32'h656c2d74 : _GEN_581;
  wire [31:0] _GEN_583 = 10'h247 == index ? 32'h2d6c6576 : _GEN_582;
  wire [31:0] _GEN_584 = 10'h248 == index ? 32'h68636163 : _GEN_583;
  wire [31:0] _GEN_585 = 10'h249 == index ? 32'h65720065 : _GEN_584;
  wire [31:0] _GEN_586 = 10'h24a == index ? 32'h69720067 : _GEN_585;
  wire [31:0] _GEN_587 = 10'h24b == index ? 32'h2c766373 : _GEN_586;
  wire [31:0] _GEN_588 = 10'h24c == index ? 32'h617369 : _GEN_587;
  wire [31:0] _GEN_589 = 10'h24d == index ? 32'h63736972 : _GEN_588;
  wire [31:0] _GEN_590 = 10'h24e == index ? 32'h6d702c76 : _GEN_589;
  wire [31:0] _GEN_591 = 10'h24f == index ? 32'h61726770 : _GEN_590;
  wire [31:0] _GEN_592 = 10'h250 == index ? 32'h616c756e : _GEN_591;
  wire [31:0] _GEN_593 = 10'h251 == index ? 32'h79746972 : _GEN_592;
  wire [31:0] _GEN_594 = 10'h252 == index ? 32'h73697200 : _GEN_593;
  wire [31:0] _GEN_595 = 10'h253 == index ? 32'h702c7663 : _GEN_594;
  wire [31:0] _GEN_596 = 10'h254 == index ? 32'h6572706d : _GEN_595;
  wire [31:0] _GEN_597 = 10'h255 == index ? 32'h6e6f6967 : _GEN_596;
  wire [31:0] _GEN_598 = 10'h256 == index ? 32'h74730073 : _GEN_597;
  wire [31:0] _GEN_599 = 10'h257 == index ? 32'h73757461 : _GEN_598;
  wire [31:0] _GEN_600 = 10'h258 == index ? 32'h626c7400 : _GEN_599;
  wire [31:0] _GEN_601 = 10'h259 == index ? 32'h6c70732d : _GEN_600;
  wire [31:0] _GEN_602 = 10'h25a == index ? 32'h23007469 : _GEN_601;
  wire [31:0] _GEN_603 = 10'h25b == index ? 32'h65746e69 : _GEN_602;
  wire [31:0] _GEN_604 = 10'h25c == index ? 32'h70757272 : _GEN_603;
  wire [31:0] _GEN_605 = 10'h25d == index ? 32'h65632d74 : _GEN_604;
  wire [31:0] _GEN_606 = 10'h25e == index ? 32'h736c6c : _GEN_605;
  wire [31:0] _GEN_607 = 10'h25f == index ? 32'h65746e69 : _GEN_606;
  wire [31:0] _GEN_608 = 10'h260 == index ? 32'h70757272 : _GEN_607;
  wire [31:0] _GEN_609 = 10'h261 == index ? 32'h6f632d74 : _GEN_608;
  wire [31:0] _GEN_610 = 10'h262 == index ? 32'h6f72746e : _GEN_609;
  wire [31:0] _GEN_611 = 10'h263 == index ? 32'h72656c6c : _GEN_610;
  wire [31:0] _GEN_612 = 10'h264 == index ? 32'h61687000 : _GEN_611;
  wire [31:0] _GEN_613 = 10'h265 == index ? 32'h656c646e : _GEN_612;
  wire [31:0] _GEN_614 = 10'h266 == index ? 32'h6e617200 : _GEN_613;
  wire [31:0] _GEN_615 = 10'h267 == index ? 32'h736567 : _GEN_614;
  wire [31:0] _GEN_616 = 10'h268 == index ? 32'h65746e69 : _GEN_615;
  wire [31:0] _GEN_617 = 10'h269 == index ? 32'h70757272 : _GEN_616;
  wire [31:0] _GEN_618 = 10'h26a == index ? 32'h652d7374 : _GEN_617;
  wire [31:0] _GEN_619 = 10'h26b == index ? 32'h6e657478 : _GEN_618;
  wire [31:0] _GEN_620 = 10'h26c == index ? 32'h646564 : _GEN_619;
  wire [31:0] _GEN_621 = 10'h26d == index ? 32'h2d676572 : _GEN_620;
  wire [31:0] _GEN_622 = 10'h26e == index ? 32'h656d616e : _GEN_621;
  wire [31:0] _GEN_623 = 10'h26f == index ? 32'h65640073 : _GEN_622;
  wire [31:0] _GEN_624 = 10'h270 == index ? 32'h2d677562 : _GEN_623;
  wire [31:0] _GEN_625 = 10'h271 == index ? 32'h61747461 : _GEN_624;
  wire [31:0] _GEN_626 = 10'h272 == index ? 32'h69006863 : _GEN_625;
  wire [31:0] _GEN_627 = 10'h273 == index ? 32'h7265746e : _GEN_626;
  wire [31:0] _GEN_628 = 10'h274 == index ? 32'h74707572 : _GEN_627;
  wire [31:0] _GEN_629 = 10'h275 == index ? 32'h7261702d : _GEN_628;
  wire [31:0] _GEN_630 = 10'h276 == index ? 32'h746e65 : _GEN_629;
  wire [31:0] _GEN_631 = 10'h277 == index ? 32'h65746e69 : _GEN_630;
  wire [31:0] _GEN_632 = 10'h278 == index ? 32'h70757272 : _GEN_631;
  wire [31:0] _GEN_633 = 10'h279 == index ? 32'h72007374 : _GEN_632;
  wire [31:0] _GEN_634 = 10'h27a == index ? 32'h76637369 : _GEN_633;
  wire [31:0] _GEN_635 = 10'h27b == index ? 32'h78616d2c : _GEN_634;
  wire [31:0] _GEN_636 = 10'h27c == index ? 32'h6972702d : _GEN_635;
  wire [31:0] _GEN_637 = 10'h27d == index ? 32'h7469726f : _GEN_636;
  wire [31:0] _GEN_638 = 10'h27e == index ? 32'h69720079 : _GEN_637;
  wire [31:0] _GEN_639 = 10'h27f == index ? 32'h2c766373 : _GEN_638;
  wire [31:0] _GEN_640 = 10'h280 == index ? 32'h7665646e : _GEN_639;
  wire [31:0] _GEN_641 = 10'h281 == index ? 32'h6c632300 : _GEN_640;
  wire [31:0] _GEN_642 = 10'h282 == index ? 32'h2d6b636f : _GEN_641;
  wire [31:0] _GEN_643 = 10'h283 == index ? 32'h6c6c6563 : _GEN_642;
  wire [31:0] _GEN_644 = 10'h284 == index ? 32'h6c630073 : _GEN_643;
  wire [31:0] _GEN_645 = 10'h285 == index ? 32'h2d6b636f : _GEN_644;
  wire [31:0] _GEN_646 = 10'h286 == index ? 32'h7074756f : _GEN_645;
  wire [31:0] _GEN_647 = 10'h287 == index ? 32'h6e2d7475 : _GEN_646;
  wire [31:0] _GEN_648 = 10'h288 == index ? 32'h73656d61 : _GEN_647;
  wire [31:0] _GEN_649 = 10'h289 == index ? 32'h0 : _GEN_648;
  wire [31:0] _GEN_650 = 10'h28a == index ? 32'h0 : _GEN_649;
  wire [31:0] _GEN_651 = 10'h28b == index ? 32'h0 : _GEN_650;
  wire [31:0] _GEN_652 = 10'h28c == index ? 32'h0 : _GEN_651;
  wire [31:0] _GEN_653 = 10'h28d == index ? 32'h0 : _GEN_652;
  wire [31:0] _GEN_654 = 10'h28e == index ? 32'h0 : _GEN_653;
  wire [31:0] _GEN_655 = 10'h28f == index ? 32'h0 : _GEN_654;
  wire [31:0] _GEN_656 = 10'h290 == index ? 32'h0 : _GEN_655;
  wire [31:0] _GEN_657 = 10'h291 == index ? 32'h0 : _GEN_656;
  wire [31:0] _GEN_658 = 10'h292 == index ? 32'h0 : _GEN_657;
  wire [31:0] _GEN_659 = 10'h293 == index ? 32'h0 : _GEN_658;
  wire [31:0] _GEN_660 = 10'h294 == index ? 32'h0 : _GEN_659;
  wire [31:0] _GEN_661 = 10'h295 == index ? 32'h0 : _GEN_660;
  wire [31:0] _GEN_662 = 10'h296 == index ? 32'h0 : _GEN_661;
  wire [31:0] _GEN_663 = 10'h297 == index ? 32'h0 : _GEN_662;
  wire [31:0] _GEN_664 = 10'h298 == index ? 32'h0 : _GEN_663;
  wire [31:0] _GEN_665 = 10'h299 == index ? 32'h0 : _GEN_664;
  wire [31:0] _GEN_666 = 10'h29a == index ? 32'h0 : _GEN_665;
  wire [31:0] _GEN_667 = 10'h29b == index ? 32'h0 : _GEN_666;
  wire [31:0] _GEN_668 = 10'h29c == index ? 32'h0 : _GEN_667;
  wire [31:0] _GEN_669 = 10'h29d == index ? 32'h0 : _GEN_668;
  wire [31:0] _GEN_670 = 10'h29e == index ? 32'h0 : _GEN_669;
  wire [31:0] _GEN_671 = 10'h29f == index ? 32'h0 : _GEN_670;
  wire [31:0] _GEN_672 = 10'h2a0 == index ? 32'h0 : _GEN_671;
  wire [31:0] _GEN_673 = 10'h2a1 == index ? 32'h0 : _GEN_672;
  wire [31:0] _GEN_674 = 10'h2a2 == index ? 32'h0 : _GEN_673;
  wire [31:0] _GEN_675 = 10'h2a3 == index ? 32'h0 : _GEN_674;
  wire [31:0] _GEN_676 = 10'h2a4 == index ? 32'h0 : _GEN_675;
  wire [31:0] _GEN_677 = 10'h2a5 == index ? 32'h0 : _GEN_676;
  wire [31:0] _GEN_678 = 10'h2a6 == index ? 32'h0 : _GEN_677;
  wire [31:0] _GEN_679 = 10'h2a7 == index ? 32'h0 : _GEN_678;
  wire [31:0] _GEN_680 = 10'h2a8 == index ? 32'h0 : _GEN_679;
  wire [31:0] _GEN_681 = 10'h2a9 == index ? 32'h0 : _GEN_680;
  wire [31:0] _GEN_682 = 10'h2aa == index ? 32'h0 : _GEN_681;
  wire [31:0] _GEN_683 = 10'h2ab == index ? 32'h0 : _GEN_682;
  wire [31:0] _GEN_684 = 10'h2ac == index ? 32'h0 : _GEN_683;
  wire [31:0] _GEN_685 = 10'h2ad == index ? 32'h0 : _GEN_684;
  wire [31:0] _GEN_686 = 10'h2ae == index ? 32'h0 : _GEN_685;
  wire [31:0] _GEN_687 = 10'h2af == index ? 32'h0 : _GEN_686;
  wire [31:0] _GEN_688 = 10'h2b0 == index ? 32'h0 : _GEN_687;
  wire [31:0] _GEN_689 = 10'h2b1 == index ? 32'h0 : _GEN_688;
  wire [31:0] _GEN_690 = 10'h2b2 == index ? 32'h0 : _GEN_689;
  wire [31:0] _GEN_691 = 10'h2b3 == index ? 32'h0 : _GEN_690;
  wire [31:0] _GEN_692 = 10'h2b4 == index ? 32'h0 : _GEN_691;
  wire [31:0] _GEN_693 = 10'h2b5 == index ? 32'h0 : _GEN_692;
  wire [31:0] _GEN_694 = 10'h2b6 == index ? 32'h0 : _GEN_693;
  wire [31:0] _GEN_695 = 10'h2b7 == index ? 32'h0 : _GEN_694;
  wire [31:0] _GEN_696 = 10'h2b8 == index ? 32'h0 : _GEN_695;
  wire [31:0] _GEN_697 = 10'h2b9 == index ? 32'h0 : _GEN_696;
  wire [31:0] _GEN_698 = 10'h2ba == index ? 32'h0 : _GEN_697;
  wire [31:0] _GEN_699 = 10'h2bb == index ? 32'h0 : _GEN_698;
  wire [31:0] _GEN_700 = 10'h2bc == index ? 32'h0 : _GEN_699;
  wire [31:0] _GEN_701 = 10'h2bd == index ? 32'h0 : _GEN_700;
  wire [31:0] _GEN_702 = 10'h2be == index ? 32'h0 : _GEN_701;
  wire [31:0] _GEN_703 = 10'h2bf == index ? 32'h0 : _GEN_702;
  wire [31:0] _GEN_704 = 10'h2c0 == index ? 32'h0 : _GEN_703;
  wire [31:0] _GEN_705 = 10'h2c1 == index ? 32'h0 : _GEN_704;
  wire [31:0] _GEN_706 = 10'h2c2 == index ? 32'h0 : _GEN_705;
  wire [31:0] _GEN_707 = 10'h2c3 == index ? 32'h0 : _GEN_706;
  wire [31:0] _GEN_708 = 10'h2c4 == index ? 32'h0 : _GEN_707;
  wire [31:0] _GEN_709 = 10'h2c5 == index ? 32'h0 : _GEN_708;
  wire [31:0] _GEN_710 = 10'h2c6 == index ? 32'h0 : _GEN_709;
  wire [31:0] _GEN_711 = 10'h2c7 == index ? 32'h0 : _GEN_710;
  wire [31:0] _GEN_712 = 10'h2c8 == index ? 32'h0 : _GEN_711;
  wire [31:0] _GEN_713 = 10'h2c9 == index ? 32'h0 : _GEN_712;
  wire [31:0] _GEN_714 = 10'h2ca == index ? 32'h0 : _GEN_713;
  wire [31:0] _GEN_715 = 10'h2cb == index ? 32'h0 : _GEN_714;
  wire [31:0] _GEN_716 = 10'h2cc == index ? 32'h0 : _GEN_715;
  wire [31:0] _GEN_717 = 10'h2cd == index ? 32'h0 : _GEN_716;
  wire [31:0] _GEN_718 = 10'h2ce == index ? 32'h0 : _GEN_717;
  wire [31:0] _GEN_719 = 10'h2cf == index ? 32'h0 : _GEN_718;
  wire [31:0] _GEN_720 = 10'h2d0 == index ? 32'h0 : _GEN_719;
  wire [31:0] _GEN_721 = 10'h2d1 == index ? 32'h0 : _GEN_720;
  wire [31:0] _GEN_722 = 10'h2d2 == index ? 32'h0 : _GEN_721;
  wire [31:0] _GEN_723 = 10'h2d3 == index ? 32'h0 : _GEN_722;
  wire [31:0] _GEN_724 = 10'h2d4 == index ? 32'h0 : _GEN_723;
  wire [31:0] _GEN_725 = 10'h2d5 == index ? 32'h0 : _GEN_724;
  wire [31:0] _GEN_726 = 10'h2d6 == index ? 32'h0 : _GEN_725;
  wire [31:0] _GEN_727 = 10'h2d7 == index ? 32'h0 : _GEN_726;
  wire [31:0] _GEN_728 = 10'h2d8 == index ? 32'h0 : _GEN_727;
  wire [31:0] _GEN_729 = 10'h2d9 == index ? 32'h0 : _GEN_728;
  wire [31:0] _GEN_730 = 10'h2da == index ? 32'h0 : _GEN_729;
  wire [31:0] _GEN_731 = 10'h2db == index ? 32'h0 : _GEN_730;
  wire [31:0] _GEN_732 = 10'h2dc == index ? 32'h0 : _GEN_731;
  wire [31:0] _GEN_733 = 10'h2dd == index ? 32'h0 : _GEN_732;
  wire [31:0] _GEN_734 = 10'h2de == index ? 32'h0 : _GEN_733;
  wire [31:0] _GEN_735 = 10'h2df == index ? 32'h0 : _GEN_734;
  wire [31:0] _GEN_736 = 10'h2e0 == index ? 32'h0 : _GEN_735;
  wire [31:0] _GEN_737 = 10'h2e1 == index ? 32'h0 : _GEN_736;
  wire [31:0] _GEN_738 = 10'h2e2 == index ? 32'h0 : _GEN_737;
  wire [31:0] _GEN_739 = 10'h2e3 == index ? 32'h0 : _GEN_738;
  wire [31:0] _GEN_740 = 10'h2e4 == index ? 32'h0 : _GEN_739;
  wire [31:0] _GEN_741 = 10'h2e5 == index ? 32'h0 : _GEN_740;
  wire [31:0] _GEN_742 = 10'h2e6 == index ? 32'h0 : _GEN_741;
  wire [31:0] _GEN_743 = 10'h2e7 == index ? 32'h0 : _GEN_742;
  wire [31:0] _GEN_744 = 10'h2e8 == index ? 32'h0 : _GEN_743;
  wire [31:0] _GEN_745 = 10'h2e9 == index ? 32'h0 : _GEN_744;
  wire [31:0] _GEN_746 = 10'h2ea == index ? 32'h0 : _GEN_745;
  wire [31:0] _GEN_747 = 10'h2eb == index ? 32'h0 : _GEN_746;
  wire [31:0] _GEN_748 = 10'h2ec == index ? 32'h0 : _GEN_747;
  wire [31:0] _GEN_749 = 10'h2ed == index ? 32'h0 : _GEN_748;
  wire [31:0] _GEN_750 = 10'h2ee == index ? 32'h0 : _GEN_749;
  wire [31:0] _GEN_751 = 10'h2ef == index ? 32'h0 : _GEN_750;
  wire [31:0] _GEN_752 = 10'h2f0 == index ? 32'h0 : _GEN_751;
  wire [31:0] _GEN_753 = 10'h2f1 == index ? 32'h0 : _GEN_752;
  wire [31:0] _GEN_754 = 10'h2f2 == index ? 32'h0 : _GEN_753;
  wire [31:0] _GEN_755 = 10'h2f3 == index ? 32'h0 : _GEN_754;
  wire [31:0] _GEN_756 = 10'h2f4 == index ? 32'h0 : _GEN_755;
  wire [31:0] _GEN_757 = 10'h2f5 == index ? 32'h0 : _GEN_756;
  wire [31:0] _GEN_758 = 10'h2f6 == index ? 32'h0 : _GEN_757;
  wire [31:0] _GEN_759 = 10'h2f7 == index ? 32'h0 : _GEN_758;
  wire [31:0] _GEN_760 = 10'h2f8 == index ? 32'h0 : _GEN_759;
  wire [31:0] _GEN_761 = 10'h2f9 == index ? 32'h0 : _GEN_760;
  wire [31:0] _GEN_762 = 10'h2fa == index ? 32'h0 : _GEN_761;
  wire [31:0] _GEN_763 = 10'h2fb == index ? 32'h0 : _GEN_762;
  wire [31:0] _GEN_764 = 10'h2fc == index ? 32'h0 : _GEN_763;
  wire [31:0] _GEN_765 = 10'h2fd == index ? 32'h0 : _GEN_764;
  wire [31:0] _GEN_766 = 10'h2fe == index ? 32'h0 : _GEN_765;
  wire [31:0] _GEN_767 = 10'h2ff == index ? 32'h0 : _GEN_766;
  wire [31:0] _GEN_768 = 10'h300 == index ? 32'h0 : _GEN_767;
  wire [31:0] _GEN_769 = 10'h301 == index ? 32'h0 : _GEN_768;
  wire [31:0] _GEN_770 = 10'h302 == index ? 32'h0 : _GEN_769;
  wire [31:0] _GEN_771 = 10'h303 == index ? 32'h0 : _GEN_770;
  wire [31:0] _GEN_772 = 10'h304 == index ? 32'h0 : _GEN_771;
  wire [31:0] _GEN_773 = 10'h305 == index ? 32'h0 : _GEN_772;
  wire [31:0] _GEN_774 = 10'h306 == index ? 32'h0 : _GEN_773;
  wire [31:0] _GEN_775 = 10'h307 == index ? 32'h0 : _GEN_774;
  wire [31:0] _GEN_776 = 10'h308 == index ? 32'h0 : _GEN_775;
  wire [31:0] _GEN_777 = 10'h309 == index ? 32'h0 : _GEN_776;
  wire [31:0] _GEN_778 = 10'h30a == index ? 32'h0 : _GEN_777;
  wire [31:0] _GEN_779 = 10'h30b == index ? 32'h0 : _GEN_778;
  wire [31:0] _GEN_780 = 10'h30c == index ? 32'h0 : _GEN_779;
  wire [31:0] _GEN_781 = 10'h30d == index ? 32'h0 : _GEN_780;
  wire [31:0] _GEN_782 = 10'h30e == index ? 32'h0 : _GEN_781;
  wire [31:0] _GEN_783 = 10'h30f == index ? 32'h0 : _GEN_782;
  wire [31:0] _GEN_784 = 10'h310 == index ? 32'h0 : _GEN_783;
  wire [31:0] _GEN_785 = 10'h311 == index ? 32'h0 : _GEN_784;
  wire [31:0] _GEN_786 = 10'h312 == index ? 32'h0 : _GEN_785;
  wire [31:0] _GEN_787 = 10'h313 == index ? 32'h0 : _GEN_786;
  wire [31:0] _GEN_788 = 10'h314 == index ? 32'h0 : _GEN_787;
  wire [31:0] _GEN_789 = 10'h315 == index ? 32'h0 : _GEN_788;
  wire [31:0] _GEN_790 = 10'h316 == index ? 32'h0 : _GEN_789;
  wire [31:0] _GEN_791 = 10'h317 == index ? 32'h0 : _GEN_790;
  wire [31:0] _GEN_792 = 10'h318 == index ? 32'h0 : _GEN_791;
  wire [31:0] _GEN_793 = 10'h319 == index ? 32'h0 : _GEN_792;
  wire [31:0] _GEN_794 = 10'h31a == index ? 32'h0 : _GEN_793;
  wire [31:0] _GEN_795 = 10'h31b == index ? 32'h0 : _GEN_794;
  wire [31:0] _GEN_796 = 10'h31c == index ? 32'h0 : _GEN_795;
  wire [31:0] _GEN_797 = 10'h31d == index ? 32'h0 : _GEN_796;
  wire [31:0] _GEN_798 = 10'h31e == index ? 32'h0 : _GEN_797;
  wire [31:0] _GEN_799 = 10'h31f == index ? 32'h0 : _GEN_798;
  wire [31:0] _GEN_800 = 10'h320 == index ? 32'h0 : _GEN_799;
  wire [31:0] _GEN_801 = 10'h321 == index ? 32'h0 : _GEN_800;
  wire [31:0] _GEN_802 = 10'h322 == index ? 32'h0 : _GEN_801;
  wire [31:0] _GEN_803 = 10'h323 == index ? 32'h0 : _GEN_802;
  wire [31:0] _GEN_804 = 10'h324 == index ? 32'h0 : _GEN_803;
  wire [31:0] _GEN_805 = 10'h325 == index ? 32'h0 : _GEN_804;
  wire [31:0] _GEN_806 = 10'h326 == index ? 32'h0 : _GEN_805;
  wire [31:0] _GEN_807 = 10'h327 == index ? 32'h0 : _GEN_806;
  wire [31:0] _GEN_808 = 10'h328 == index ? 32'h0 : _GEN_807;
  wire [31:0] _GEN_809 = 10'h329 == index ? 32'h0 : _GEN_808;
  wire [31:0] _GEN_810 = 10'h32a == index ? 32'h0 : _GEN_809;
  wire [31:0] _GEN_811 = 10'h32b == index ? 32'h0 : _GEN_810;
  wire [31:0] _GEN_812 = 10'h32c == index ? 32'h0 : _GEN_811;
  wire [31:0] _GEN_813 = 10'h32d == index ? 32'h0 : _GEN_812;
  wire [31:0] _GEN_814 = 10'h32e == index ? 32'h0 : _GEN_813;
  wire [31:0] _GEN_815 = 10'h32f == index ? 32'h0 : _GEN_814;
  wire [31:0] _GEN_816 = 10'h330 == index ? 32'h0 : _GEN_815;
  wire [31:0] _GEN_817 = 10'h331 == index ? 32'h0 : _GEN_816;
  wire [31:0] _GEN_818 = 10'h332 == index ? 32'h0 : _GEN_817;
  wire [31:0] _GEN_819 = 10'h333 == index ? 32'h0 : _GEN_818;
  wire [31:0] _GEN_820 = 10'h334 == index ? 32'h0 : _GEN_819;
  wire [31:0] _GEN_821 = 10'h335 == index ? 32'h0 : _GEN_820;
  wire [31:0] _GEN_822 = 10'h336 == index ? 32'h0 : _GEN_821;
  wire [31:0] _GEN_823 = 10'h337 == index ? 32'h0 : _GEN_822;
  wire [31:0] _GEN_824 = 10'h338 == index ? 32'h0 : _GEN_823;
  wire [31:0] _GEN_825 = 10'h339 == index ? 32'h0 : _GEN_824;
  wire [31:0] _GEN_826 = 10'h33a == index ? 32'h0 : _GEN_825;
  wire [31:0] _GEN_827 = 10'h33b == index ? 32'h0 : _GEN_826;
  wire [31:0] _GEN_828 = 10'h33c == index ? 32'h0 : _GEN_827;
  wire [31:0] _GEN_829 = 10'h33d == index ? 32'h0 : _GEN_828;
  wire [31:0] _GEN_830 = 10'h33e == index ? 32'h0 : _GEN_829;
  wire [31:0] _GEN_831 = 10'h33f == index ? 32'h0 : _GEN_830;
  wire [31:0] _GEN_832 = 10'h340 == index ? 32'h0 : _GEN_831;
  wire [31:0] _GEN_833 = 10'h341 == index ? 32'h0 : _GEN_832;
  wire [31:0] _GEN_834 = 10'h342 == index ? 32'h0 : _GEN_833;
  wire [31:0] _GEN_835 = 10'h343 == index ? 32'h0 : _GEN_834;
  wire [31:0] _GEN_836 = 10'h344 == index ? 32'h0 : _GEN_835;
  wire [31:0] _GEN_837 = 10'h345 == index ? 32'h0 : _GEN_836;
  wire [31:0] _GEN_838 = 10'h346 == index ? 32'h0 : _GEN_837;
  wire [31:0] _GEN_839 = 10'h347 == index ? 32'h0 : _GEN_838;
  wire [31:0] _GEN_840 = 10'h348 == index ? 32'h0 : _GEN_839;
  wire [31:0] _GEN_841 = 10'h349 == index ? 32'h0 : _GEN_840;
  wire [31:0] _GEN_842 = 10'h34a == index ? 32'h0 : _GEN_841;
  wire [31:0] _GEN_843 = 10'h34b == index ? 32'h0 : _GEN_842;
  wire [31:0] _GEN_844 = 10'h34c == index ? 32'h0 : _GEN_843;
  wire [31:0] _GEN_845 = 10'h34d == index ? 32'h0 : _GEN_844;
  wire [31:0] _GEN_846 = 10'h34e == index ? 32'h0 : _GEN_845;
  wire [31:0] _GEN_847 = 10'h34f == index ? 32'h0 : _GEN_846;
  wire [31:0] _GEN_848 = 10'h350 == index ? 32'h0 : _GEN_847;
  wire [31:0] _GEN_849 = 10'h351 == index ? 32'h0 : _GEN_848;
  wire [31:0] _GEN_850 = 10'h352 == index ? 32'h0 : _GEN_849;
  wire [31:0] _GEN_851 = 10'h353 == index ? 32'h0 : _GEN_850;
  wire [31:0] _GEN_852 = 10'h354 == index ? 32'h0 : _GEN_851;
  wire [31:0] _GEN_853 = 10'h355 == index ? 32'h0 : _GEN_852;
  wire [31:0] _GEN_854 = 10'h356 == index ? 32'h0 : _GEN_853;
  wire [31:0] _GEN_855 = 10'h357 == index ? 32'h0 : _GEN_854;
  wire [31:0] _GEN_856 = 10'h358 == index ? 32'h0 : _GEN_855;
  wire [31:0] _GEN_857 = 10'h359 == index ? 32'h0 : _GEN_856;
  wire [31:0] _GEN_858 = 10'h35a == index ? 32'h0 : _GEN_857;
  wire [31:0] _GEN_859 = 10'h35b == index ? 32'h0 : _GEN_858;
  wire [31:0] _GEN_860 = 10'h35c == index ? 32'h0 : _GEN_859;
  wire [31:0] _GEN_861 = 10'h35d == index ? 32'h0 : _GEN_860;
  wire [31:0] _GEN_862 = 10'h35e == index ? 32'h0 : _GEN_861;
  wire [31:0] _GEN_863 = 10'h35f == index ? 32'h0 : _GEN_862;
  wire [31:0] _GEN_864 = 10'h360 == index ? 32'h0 : _GEN_863;
  wire [31:0] _GEN_865 = 10'h361 == index ? 32'h0 : _GEN_864;
  wire [31:0] _GEN_866 = 10'h362 == index ? 32'h0 : _GEN_865;
  wire [31:0] _GEN_867 = 10'h363 == index ? 32'h0 : _GEN_866;
  wire [31:0] _GEN_868 = 10'h364 == index ? 32'h0 : _GEN_867;
  wire [31:0] _GEN_869 = 10'h365 == index ? 32'h0 : _GEN_868;
  wire [31:0] _GEN_870 = 10'h366 == index ? 32'h0 : _GEN_869;
  wire [31:0] _GEN_871 = 10'h367 == index ? 32'h0 : _GEN_870;
  wire [31:0] _GEN_872 = 10'h368 == index ? 32'h0 : _GEN_871;
  wire [31:0] _GEN_873 = 10'h369 == index ? 32'h0 : _GEN_872;
  wire [31:0] _GEN_874 = 10'h36a == index ? 32'h0 : _GEN_873;
  wire [31:0] _GEN_875 = 10'h36b == index ? 32'h0 : _GEN_874;
  wire [31:0] _GEN_876 = 10'h36c == index ? 32'h0 : _GEN_875;
  wire [31:0] _GEN_877 = 10'h36d == index ? 32'h0 : _GEN_876;
  wire [31:0] _GEN_878 = 10'h36e == index ? 32'h0 : _GEN_877;
  wire [31:0] _GEN_879 = 10'h36f == index ? 32'h0 : _GEN_878;
  wire [31:0] _GEN_880 = 10'h370 == index ? 32'h0 : _GEN_879;
  wire [31:0] _GEN_881 = 10'h371 == index ? 32'h0 : _GEN_880;
  wire [31:0] _GEN_882 = 10'h372 == index ? 32'h0 : _GEN_881;
  wire [31:0] _GEN_883 = 10'h373 == index ? 32'h0 : _GEN_882;
  wire [31:0] _GEN_884 = 10'h374 == index ? 32'h0 : _GEN_883;
  wire [31:0] _GEN_885 = 10'h375 == index ? 32'h0 : _GEN_884;
  wire [31:0] _GEN_886 = 10'h376 == index ? 32'h0 : _GEN_885;
  wire [31:0] _GEN_887 = 10'h377 == index ? 32'h0 : _GEN_886;
  wire [31:0] _GEN_888 = 10'h378 == index ? 32'h0 : _GEN_887;
  wire [31:0] _GEN_889 = 10'h379 == index ? 32'h0 : _GEN_888;
  wire [31:0] _GEN_890 = 10'h37a == index ? 32'h0 : _GEN_889;
  wire [31:0] _GEN_891 = 10'h37b == index ? 32'h0 : _GEN_890;
  wire [31:0] _GEN_892 = 10'h37c == index ? 32'h0 : _GEN_891;
  wire [31:0] _GEN_893 = 10'h37d == index ? 32'h0 : _GEN_892;
  wire [31:0] _GEN_894 = 10'h37e == index ? 32'h0 : _GEN_893;
  wire [31:0] _GEN_895 = 10'h37f == index ? 32'h0 : _GEN_894;
  wire [31:0] _GEN_896 = 10'h380 == index ? 32'h0 : _GEN_895;
  wire [31:0] _GEN_897 = 10'h381 == index ? 32'h0 : _GEN_896;
  wire [31:0] _GEN_898 = 10'h382 == index ? 32'h0 : _GEN_897;
  wire [31:0] _GEN_899 = 10'h383 == index ? 32'h0 : _GEN_898;
  wire [31:0] _GEN_900 = 10'h384 == index ? 32'h0 : _GEN_899;
  wire [31:0] _GEN_901 = 10'h385 == index ? 32'h0 : _GEN_900;
  wire [31:0] _GEN_902 = 10'h386 == index ? 32'h0 : _GEN_901;
  wire [31:0] _GEN_903 = 10'h387 == index ? 32'h0 : _GEN_902;
  wire [31:0] _GEN_904 = 10'h388 == index ? 32'h0 : _GEN_903;
  wire [31:0] _GEN_905 = 10'h389 == index ? 32'h0 : _GEN_904;
  wire [31:0] _GEN_906 = 10'h38a == index ? 32'h0 : _GEN_905;
  wire [31:0] _GEN_907 = 10'h38b == index ? 32'h0 : _GEN_906;
  wire [31:0] _GEN_908 = 10'h38c == index ? 32'h0 : _GEN_907;
  wire [31:0] _GEN_909 = 10'h38d == index ? 32'h0 : _GEN_908;
  wire [31:0] _GEN_910 = 10'h38e == index ? 32'h0 : _GEN_909;
  wire [31:0] _GEN_911 = 10'h38f == index ? 32'h0 : _GEN_910;
  wire [31:0] _GEN_912 = 10'h390 == index ? 32'h0 : _GEN_911;
  wire [31:0] _GEN_913 = 10'h391 == index ? 32'h0 : _GEN_912;
  wire [31:0] _GEN_914 = 10'h392 == index ? 32'h0 : _GEN_913;
  wire [31:0] _GEN_915 = 10'h393 == index ? 32'h0 : _GEN_914;
  wire [31:0] _GEN_916 = 10'h394 == index ? 32'h0 : _GEN_915;
  wire [31:0] _GEN_917 = 10'h395 == index ? 32'h0 : _GEN_916;
  wire [31:0] _GEN_918 = 10'h396 == index ? 32'h0 : _GEN_917;
  wire [31:0] _GEN_919 = 10'h397 == index ? 32'h0 : _GEN_918;
  wire [31:0] _GEN_920 = 10'h398 == index ? 32'h0 : _GEN_919;
  wire [31:0] _GEN_921 = 10'h399 == index ? 32'h0 : _GEN_920;
  wire [31:0] _GEN_922 = 10'h39a == index ? 32'h0 : _GEN_921;
  wire [31:0] _GEN_923 = 10'h39b == index ? 32'h0 : _GEN_922;
  wire [31:0] _GEN_924 = 10'h39c == index ? 32'h0 : _GEN_923;
  wire [31:0] _GEN_925 = 10'h39d == index ? 32'h0 : _GEN_924;
  wire [31:0] _GEN_926 = 10'h39e == index ? 32'h0 : _GEN_925;
  wire [31:0] _GEN_927 = 10'h39f == index ? 32'h0 : _GEN_926;
  wire [31:0] _GEN_928 = 10'h3a0 == index ? 32'h0 : _GEN_927;
  wire [31:0] _GEN_929 = 10'h3a1 == index ? 32'h0 : _GEN_928;
  wire [31:0] _GEN_930 = 10'h3a2 == index ? 32'h0 : _GEN_929;
  wire [31:0] _GEN_931 = 10'h3a3 == index ? 32'h0 : _GEN_930;
  wire [31:0] _GEN_932 = 10'h3a4 == index ? 32'h0 : _GEN_931;
  wire [31:0] _GEN_933 = 10'h3a5 == index ? 32'h0 : _GEN_932;
  wire [31:0] _GEN_934 = 10'h3a6 == index ? 32'h0 : _GEN_933;
  wire [31:0] _GEN_935 = 10'h3a7 == index ? 32'h0 : _GEN_934;
  wire [31:0] _GEN_936 = 10'h3a8 == index ? 32'h0 : _GEN_935;
  wire [31:0] _GEN_937 = 10'h3a9 == index ? 32'h0 : _GEN_936;
  wire [31:0] _GEN_938 = 10'h3aa == index ? 32'h0 : _GEN_937;
  wire [31:0] _GEN_939 = 10'h3ab == index ? 32'h0 : _GEN_938;
  wire [31:0] _GEN_940 = 10'h3ac == index ? 32'h0 : _GEN_939;
  wire [31:0] _GEN_941 = 10'h3ad == index ? 32'h0 : _GEN_940;
  wire [31:0] _GEN_942 = 10'h3ae == index ? 32'h0 : _GEN_941;
  wire [31:0] _GEN_943 = 10'h3af == index ? 32'h0 : _GEN_942;
  wire [31:0] _GEN_944 = 10'h3b0 == index ? 32'h0 : _GEN_943;
  wire [31:0] _GEN_945 = 10'h3b1 == index ? 32'h0 : _GEN_944;
  wire [31:0] _GEN_946 = 10'h3b2 == index ? 32'h0 : _GEN_945;
  wire [31:0] _GEN_947 = 10'h3b3 == index ? 32'h0 : _GEN_946;
  wire [31:0] _GEN_948 = 10'h3b4 == index ? 32'h0 : _GEN_947;
  wire [31:0] _GEN_949 = 10'h3b5 == index ? 32'h0 : _GEN_948;
  wire [31:0] _GEN_950 = 10'h3b6 == index ? 32'h0 : _GEN_949;
  wire [31:0] _GEN_951 = 10'h3b7 == index ? 32'h0 : _GEN_950;
  wire [31:0] _GEN_952 = 10'h3b8 == index ? 32'h0 : _GEN_951;
  wire [31:0] _GEN_953 = 10'h3b9 == index ? 32'h0 : _GEN_952;
  wire [31:0] _GEN_954 = 10'h3ba == index ? 32'h0 : _GEN_953;
  wire [31:0] _GEN_955 = 10'h3bb == index ? 32'h0 : _GEN_954;
  wire [31:0] _GEN_956 = 10'h3bc == index ? 32'h0 : _GEN_955;
  wire [31:0] _GEN_957 = 10'h3bd == index ? 32'h0 : _GEN_956;
  wire [31:0] _GEN_958 = 10'h3be == index ? 32'h0 : _GEN_957;
  wire [31:0] _GEN_959 = 10'h3bf == index ? 32'h0 : _GEN_958;
  wire [31:0] _GEN_960 = 10'h3c0 == index ? 32'h0 : _GEN_959;
  wire [31:0] _GEN_961 = 10'h3c1 == index ? 32'h0 : _GEN_960;
  wire [31:0] _GEN_962 = 10'h3c2 == index ? 32'h0 : _GEN_961;
  wire [31:0] _GEN_963 = 10'h3c3 == index ? 32'h0 : _GEN_962;
  wire [31:0] _GEN_964 = 10'h3c4 == index ? 32'h0 : _GEN_963;
  wire [31:0] _GEN_965 = 10'h3c5 == index ? 32'h0 : _GEN_964;
  wire [31:0] _GEN_966 = 10'h3c6 == index ? 32'h0 : _GEN_965;
  wire [31:0] _GEN_967 = 10'h3c7 == index ? 32'h0 : _GEN_966;
  wire [31:0] _GEN_968 = 10'h3c8 == index ? 32'h0 : _GEN_967;
  wire [31:0] _GEN_969 = 10'h3c9 == index ? 32'h0 : _GEN_968;
  wire [31:0] _GEN_970 = 10'h3ca == index ? 32'h0 : _GEN_969;
  wire [31:0] _GEN_971 = 10'h3cb == index ? 32'h0 : _GEN_970;
  wire [31:0] _GEN_972 = 10'h3cc == index ? 32'h0 : _GEN_971;
  wire [31:0] _GEN_973 = 10'h3cd == index ? 32'h0 : _GEN_972;
  wire [31:0] _GEN_974 = 10'h3ce == index ? 32'h0 : _GEN_973;
  wire [31:0] _GEN_975 = 10'h3cf == index ? 32'h0 : _GEN_974;
  wire [31:0] _GEN_976 = 10'h3d0 == index ? 32'h0 : _GEN_975;
  wire [31:0] _GEN_977 = 10'h3d1 == index ? 32'h0 : _GEN_976;
  wire [31:0] _GEN_978 = 10'h3d2 == index ? 32'h0 : _GEN_977;
  wire [31:0] _GEN_979 = 10'h3d3 == index ? 32'h0 : _GEN_978;
  wire [31:0] _GEN_980 = 10'h3d4 == index ? 32'h0 : _GEN_979;
  wire [31:0] _GEN_981 = 10'h3d5 == index ? 32'h0 : _GEN_980;
  wire [31:0] _GEN_982 = 10'h3d6 == index ? 32'h0 : _GEN_981;
  wire [31:0] _GEN_983 = 10'h3d7 == index ? 32'h0 : _GEN_982;
  wire [31:0] _GEN_984 = 10'h3d8 == index ? 32'h0 : _GEN_983;
  wire [31:0] _GEN_985 = 10'h3d9 == index ? 32'h0 : _GEN_984;
  wire [31:0] _GEN_986 = 10'h3da == index ? 32'h0 : _GEN_985;
  wire [31:0] _GEN_987 = 10'h3db == index ? 32'h0 : _GEN_986;
  wire [31:0] _GEN_988 = 10'h3dc == index ? 32'h0 : _GEN_987;
  wire [31:0] _GEN_989 = 10'h3dd == index ? 32'h0 : _GEN_988;
  wire [31:0] _GEN_990 = 10'h3de == index ? 32'h0 : _GEN_989;
  wire [31:0] _GEN_991 = 10'h3df == index ? 32'h0 : _GEN_990;
  wire [31:0] _GEN_992 = 10'h3e0 == index ? 32'h0 : _GEN_991;
  wire [31:0] _GEN_993 = 10'h3e1 == index ? 32'h0 : _GEN_992;
  wire [31:0] _GEN_994 = 10'h3e2 == index ? 32'h0 : _GEN_993;
  wire [31:0] _GEN_995 = 10'h3e3 == index ? 32'h0 : _GEN_994;
  wire [31:0] _GEN_996 = 10'h3e4 == index ? 32'h0 : _GEN_995;
  wire [31:0] _GEN_997 = 10'h3e5 == index ? 32'h0 : _GEN_996;
  wire [31:0] _GEN_998 = 10'h3e6 == index ? 32'h0 : _GEN_997;
  wire [31:0] _GEN_999 = 10'h3e7 == index ? 32'h0 : _GEN_998;
  wire [31:0] _GEN_1000 = 10'h3e8 == index ? 32'h0 : _GEN_999;
  wire [31:0] _GEN_1001 = 10'h3e9 == index ? 32'h0 : _GEN_1000;
  wire [31:0] _GEN_1002 = 10'h3ea == index ? 32'h0 : _GEN_1001;
  wire [31:0] _GEN_1003 = 10'h3eb == index ? 32'h0 : _GEN_1002;
  wire [31:0] _GEN_1004 = 10'h3ec == index ? 32'h0 : _GEN_1003;
  wire [31:0] _GEN_1005 = 10'h3ed == index ? 32'h0 : _GEN_1004;
  wire [31:0] _GEN_1006 = 10'h3ee == index ? 32'h0 : _GEN_1005;
  wire [31:0] _GEN_1007 = 10'h3ef == index ? 32'h0 : _GEN_1006;
  wire [31:0] _GEN_1008 = 10'h3f0 == index ? 32'h0 : _GEN_1007;
  wire [31:0] _GEN_1009 = 10'h3f1 == index ? 32'h0 : _GEN_1008;
  wire [31:0] _GEN_1010 = 10'h3f2 == index ? 32'h0 : _GEN_1009;
  wire [31:0] _GEN_1011 = 10'h3f3 == index ? 32'h0 : _GEN_1010;
  wire [31:0] _GEN_1012 = 10'h3f4 == index ? 32'h0 : _GEN_1011;
  wire [31:0] _GEN_1013 = 10'h3f5 == index ? 32'h0 : _GEN_1012;
  wire [31:0] _GEN_1014 = 10'h3f6 == index ? 32'h0 : _GEN_1013;
  wire [31:0] _GEN_1015 = 10'h3f7 == index ? 32'h0 : _GEN_1014;
  wire [31:0] _GEN_1016 = 10'h3f8 == index ? 32'h0 : _GEN_1015;
  wire [31:0] _GEN_1017 = 10'h3f9 == index ? 32'h0 : _GEN_1016;
  wire [31:0] _GEN_1018 = 10'h3fa == index ? 32'h0 : _GEN_1017;
  wire [31:0] _GEN_1019 = 10'h3fb == index ? 32'h0 : _GEN_1018;
  wire [31:0] _GEN_1020 = 10'h3fc == index ? 32'h0 : _GEN_1019;
  wire [31:0] _GEN_1021 = 10'h3fd == index ? 32'h0 : _GEN_1020;
  wire [31:0] _GEN_1022 = 10'h3fe == index ? 32'h0 : _GEN_1021;
  wire [31:0] _GEN_1023 = 10'h3ff == index ? 32'h0 : _GEN_1022;
  
  assign auto_in_a_ready = auto_in_d_ready;
  assign auto_in_d_valid = auto_in_a_valid;
  assign auto_in_d_bits_size = auto_in_a_bits_size;
  assign auto_in_d_bits_source = auto_in_a_bits_source;
  assign auto_in_d_bits_data = |high ? 32'h0 : _GEN_1023;
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = auto_in_d_ready;
  assign monitor_io_in_a_valid = auto_in_a_valid;
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
  assign monitor_io_in_d_ready = auto_in_d_ready;
  assign monitor_io_in_d_valid = auto_in_a_valid;
  assign monitor_io_in_d_bits_size = auto_in_a_bits_size;
  assign monitor_io_in_d_bits_source = auto_in_a_bits_source;
endmodule