// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`default_nettype wire




module RVX_MODULE_042(
  input         rvx_port_25,
  input         rvx_port_41,
  input         rvx_port_26,
  input         rvx_port_03,
  input         rvx_port_30,
  input         rvx_port_35,
  input         rvx_port_13,
  input         rvx_port_19,
  input         rvx_port_29,
  input         rvx_port_32,
  input         rvx_port_28,
  input         rvx_port_17,
  input         rvx_port_12,
  input         rvx_port_48,
  input         rvx_port_37,
  input         rvx_port_43,
  input         rvx_port_01,
  input         rvx_port_09,
  input         rvx_port_05,
  input         rvx_port_08,
  input         rvx_port_11,
  input         rvx_port_47,
  input         rvx_port_15,
  input         rvx_port_07,
  input         rvx_port_23,
  input         rvx_port_36,
  input         rvx_port_10,
  input         rvx_port_06,
  input         rvx_port_20,
  input         rvx_port_44,
  input         rvx_port_02,
  input         rvx_port_00,
  input         rvx_port_21,
  input         rvx_port_16,
  output        rvx_port_22,
  output        rvx_port_40,
  input         rvx_port_34,
  input  [2:0]  rvx_port_18,
  input  [1:0]  rvx_port_04,
  input  [9:0]  rvx_port_42,
  input  [27:0] rvx_port_45,
  input  [3:0]  rvx_port_38,
  input  [31:0] rvx_port_33,
  input         rvx_port_31,
  output        rvx_port_27,
  output [2:0]  rvx_port_39,
  output [1:0]  rvx_port_14,
  output [9:0]  rvx_port_46,
  output [31:0] rvx_port_24
);



  wire  _T_31_a_ready;
  wire  _T_31_a_valid;
  wire [2:0] _T_31_a_bits_opcode;
  wire [1:0] _T_31_a_bits_size;
  wire [9:0] _T_31_a_bits_source;
  wire [27:0] _T_31_a_bits_address;
  wire [3:0] _T_31_a_bits_mask;
  wire [31:0] _T_31_a_bits_data;
  wire  _T_31_d_ready;
  wire  _T_31_d_valid;
  wire [2:0] _T_31_d_bits_opcode;
  wire [1:0] _T_31_d_bits_size;
  wire [9:0] _T_31_d_bits_source;
  wire [31:0] _T_31_d_bits_data;
  wire  rvx_signal_455;
  wire  rvx_signal_394;
  wire  rvx_signal_082;
  wire  rvx_signal_031;
  wire  rvx_signal_112;
  wire  rvx_signal_169;
  wire  rvx_signal_288;
  wire  rvx_signal_353;
  wire  rvx_signal_216;
  wire  rvx_signal_419;
  wire  rvx_signal_109;
  wire  rvx_signal_458;
  wire  rvx_signal_411;
  wire  rvx_signal_412;
  wire  rvx_signal_262;
  wire  rvx_signal_367;
  wire  rvx_signal_200;
  wire  rvx_signal_046;
  wire  rvx_signal_403;
  wire  rvx_signal_402;
  wire  rvx_signal_193;
  wire  rvx_signal_154;
  wire  rvx_signal_325;
  wire  rvx_signal_381;
  wire  rvx_signal_348;
  wire  rvx_signal_334;
  wire  rvx_signal_102;
  wire  rvx_signal_323;
  wire  rvx_signal_231;
  wire  rvx_signal_115;
  wire  rvx_signal_218;
  wire  rvx_signal_122;
  wire  rvx_signal_448;
  wire  rvx_signal_108;
  wire  rvx_signal_006;
  wire  rvx_signal_123;
  wire  rvx_signal_259;
  wire  rvx_signal_256;
  wire  rvx_signal_130;
  wire  rvx_signal_098;
  wire  rvx_signal_081;
  wire  rvx_signal_149;
  wire  rvx_signal_307;
  wire  rvx_signal_075;
  wire  rvx_signal_027;
  wire  rvx_signal_012;
  wire  rvx_signal_327;
  wire  rvx_signal_441;
  wire  rvx_signal_146;
  wire  rvx_signal_452;
  wire  rvx_signal_428;
  wire  rvx_signal_338;
  wire  rvx_signal_203;
  wire  rvx_signal_461;
  wire  rvx_signal_152;
  wire  rvx_signal_101;
  wire  rvx_signal_244;
  wire  rvx_signal_159;
  wire  rvx_signal_054;
  wire  rvx_signal_000;
  wire  rvx_signal_321;
  wire  rvx_signal_024;
  wire  rvx_signal_174;
  wire  rvx_signal_360;
  wire  rvx_signal_297;
  wire  rvx_signal_036;
  wire  rvx_signal_100;
  wire  rvx_signal_341;
  wire  rvx_signal_209;
  wire  rvx_signal_401;
  wire  rvx_signal_425;
  wire  rvx_signal_198;
  wire  rvx_signal_285;
  wire  rvx_signal_326;
  wire  rvx_signal_201;
  wire  rvx_signal_451;
  wire  rvx_signal_074;
  wire  rvx_signal_063;
  wire  rvx_signal_087;
  wire  rvx_signal_186;
  wire  rvx_signal_379;
  wire  rvx_signal_204;
  wire  rvx_signal_405;
  wire  rvx_signal_192;
  wire  rvx_signal_366;
  wire  rvx_signal_312;
  wire  rvx_signal_282;
  wire  rvx_signal_125;
  wire  rvx_signal_330;
  wire  rvx_signal_148;
  wire  rvx_signal_195;
  wire  rvx_signal_180;
  wire  rvx_signal_295;
  wire  rvx_signal_085;
  wire  rvx_signal_163;
  wire  rvx_signal_336;
  wire  rvx_signal_449;
  wire  rvx_signal_254;
  wire  rvx_signal_391;
  wire  rvx_signal_390;
  wire  rvx_signal_439;
  wire  rvx_signal_028;
  wire  rvx_signal_363;
  wire  rvx_signal_062;
  wire  rvx_signal_220;
  wire  rvx_signal_299;
  wire  rvx_signal_128;
  wire  rvx_signal_141;
  wire  rvx_signal_143;
  wire  rvx_signal_226;
  wire  rvx_signal_347;
  wire  rvx_signal_070;
  wire  rvx_signal_039;
  wire  rvx_signal_213;
  wire  rvx_signal_056;
  wire  rvx_signal_090;
  wire  rvx_signal_151;
  wire  rvx_signal_042;
  wire  rvx_signal_464;
  wire  rvx_signal_135;
  wire  rvx_signal_083;
  wire  rvx_signal_127;
  wire  rvx_signal_206;
  wire  rvx_signal_235;
  wire  rvx_signal_156;
  wire  rvx_signal_010;
  wire  rvx_signal_314;
  wire  rvx_signal_053;
  wire  rvx_signal_252;
  wire  rvx_signal_044;
  wire  rvx_signal_398;
  wire  rvx_signal_227;
  wire  rvx_signal_283;
  wire  rvx_signal_373;
  wire  rvx_signal_041;
  wire  rvx_signal_308;
  wire  rvx_signal_463;
  wire  rvx_signal_368;
  wire  rvx_signal_345;
  wire  rvx_signal_037;
  wire  rvx_signal_356;
  wire  rvx_signal_187;
  wire  rvx_signal_317;
  wire  rvx_signal_236;
  wire  rvx_signal_292;
  wire  rvx_signal_093;
  wire  rvx_signal_471;
  wire  rvx_signal_413;
  wire  rvx_signal_013;
  wire  rvx_signal_301;
  wire  rvx_signal_136;
  wire  rvx_signal_177;
  wire  rvx_signal_324;
  wire  rvx_signal_474;
  wire  rvx_signal_107;
  wire  rvx_signal_343;
  wire  rvx_signal_328;
  wire  rvx_signal_389;
  wire  rvx_signal_337;
  wire  rvx_signal_015;
  wire  rvx_signal_095;
  wire  rvx_signal_477;
  wire  rvx_signal_188;
  wire  rvx_signal_030;
  wire  rvx_signal_459;
  wire  rvx_signal_468;
  wire  rvx_signal_084;
  wire  rvx_signal_194;
  wire  rvx_signal_132;
  wire  rvx_signal_424;
  wire  rvx_signal_329;
  wire  rvx_signal_291;
  wire  rvx_signal_051;
  wire  rvx_signal_175;
  wire  rvx_signal_406;
  wire  rvx_signal_223;
  wire  rvx_signal_205;
  wire  rvx_signal_257;
  wire  rvx_signal_361;
  wire  rvx_signal_352;
  wire  rvx_signal_466;
  wire  rvx_signal_442;
  wire  rvx_signal_335;
  wire  rvx_signal_417;
  wire  rvx_signal_217;
  wire  rvx_signal_438;
  wire  rvx_signal_014;
  wire  rvx_signal_104;
  wire  rvx_signal_219;
  wire  rvx_signal_133;
  wire  rvx_signal_142;
  wire  rvx_signal_380;
  wire  rvx_signal_344;
  wire  rvx_signal_113;
  wire  rvx_signal_310;
  wire  rvx_signal_079;
  wire  rvx_signal_049;
  wire  rvx_signal_091;
  wire  rvx_signal_208;
  wire  rvx_signal_346;
  wire  rvx_signal_246;
  wire  rvx_signal_214;
  wire  rvx_signal_261;
  wire  rvx_signal_355;
  wire  rvx_signal_278;
  wire  rvx_signal_440;
  wire  rvx_signal_157;
  wire  rvx_signal_434;
  wire  rvx_signal_293;
  wire  rvx_signal_021;
  wire  rvx_signal_268;
  wire  rvx_signal_320;
  wire  rvx_signal_076;
  wire  rvx_signal_016;
  wire  rvx_signal_281;
  wire  rvx_signal_393;
  wire  rvx_signal_168;
  wire  rvx_signal_270;
  wire  rvx_signal_376;
  wire  rvx_signal_375;
  wire  rvx_signal_362;
  wire  rvx_signal_121;
  wire  rvx_signal_196;
  wire  rvx_signal_009;
  wire  rvx_signal_237;
  wire  rvx_signal_385;
  wire  rvx_signal_331;
  wire  rvx_signal_210;
  wire  rvx_signal_271;
  wire  rvx_signal_284;
  wire  rvx_signal_073;
  wire  rvx_signal_280;
  wire  rvx_signal_269;
  wire  rvx_signal_047;
  wire  rvx_signal_158;
  wire  rvx_signal_119;
  wire  rvx_signal_414;
  wire  rvx_signal_357;
  wire  rvx_signal_184;
  wire  rvx_signal_313;
  wire  rvx_signal_055;
  wire  rvx_signal_251;
  wire  rvx_signal_170;
  wire  rvx_signal_420;
  wire  rvx_signal_199;
  wire  rvx_signal_277;
  wire  rvx_signal_453;
  wire  rvx_signal_378;
  wire  rvx_signal_040;
  wire  rvx_signal_377;
  wire  rvx_signal_349;
  wire  rvx_signal_447;
  wire  rvx_signal_106;
  wire  rvx_signal_241;
  wire  rvx_signal_078;
  wire  rvx_signal_134;
  wire  rvx_signal_365;
  wire  rvx_signal_457;
  wire  rvx_signal_138;
  wire  rvx_signal_422;
  wire  rvx_signal_472;
  wire  rvx_signal_387;
  wire  rvx_signal_351;
  wire  rvx_signal_212;
  wire  rvx_signal_069;
  wire  rvx_signal_068;
  wire  rvx_signal_473;
  wire  rvx_signal_160;
  wire  rvx_signal_118;
  wire  rvx_signal_397;
  wire  rvx_signal_035;
  wire  rvx_signal_305;
  wire  rvx_signal_340;
  wire  rvx_signal_421;
  wire  rvx_signal_233;
  wire  rvx_signal_247;
  wire  rvx_signal_333;
  wire  rvx_signal_022;
  wire  rvx_signal_274;
  wire  rvx_signal_020;
  wire  rvx_signal_086;
  wire  rvx_signal_211;
  wire  rvx_signal_207;
  wire  rvx_signal_416;
  wire  rvx_signal_171;
  wire  rvx_signal_354;
  wire  rvx_signal_190;
  wire  rvx_signal_071;
  wire  rvx_signal_392;
  wire  rvx_signal_225;
  wire  rvx_signal_094;
  wire  rvx_signal_176;
  wire  rvx_signal_469;
  wire  rvx_signal_139;
  wire  rvx_signal_264;
  wire  rvx_signal_460;
  wire  rvx_signal_191;
  wire  rvx_signal_302;
  wire  rvx_signal_404;
  wire  rvx_signal_147;
  wire  rvx_signal_342;
  wire  rvx_signal_315;
  wire  rvx_signal_105;
  wire  rvx_signal_467;
  wire  rvx_signal_003;
  wire  rvx_signal_396;
  wire  rvx_signal_250;
  wire  rvx_signal_181;
  wire  rvx_signal_059;
  wire  rvx_signal_476;
  wire  rvx_signal_287;
  wire  rvx_signal_319;
  wire  rvx_signal_026;
  wire  rvx_signal_072;
  wire  rvx_signal_260;
  wire  rvx_signal_478;
  wire  rvx_signal_276;
  wire  rvx_signal_322;
  wire  rvx_signal_230;
  wire  rvx_signal_273;
  wire  rvx_signal_456;
  wire  rvx_signal_232;
  wire  rvx_signal_445;
  wire  rvx_signal_061;
  wire  rvx_signal_370;
  wire  rvx_signal_173;
  wire  rvx_signal_286;
  wire  rvx_signal_339;
  reg [2:0] rvx_signal_243;

  reg [2:0] rvx_signal_057;

  reg [2:0] rvx_signal_311;

  reg [2:0] rvx_signal_089;

  reg [2:0] rvx_signal_117;

  reg [2:0] rvx_signal_116;

  reg [2:0] rvx_signal_415;

  reg [2:0] rvx_signal_289;

  reg [2:0] rvx_signal_002;

  reg [2:0] rvx_signal_395;

  reg [2:0] rvx_signal_140;

  reg [2:0] rvx_signal_023;

  reg [2:0] rvx_signal_145;

  reg [2:0] rvx_signal_025;

  reg [2:0] rvx_signal_418;

  reg [2:0] rvx_signal_008;

  reg [2:0] rvx_signal_245;

  reg [2:0] rvx_signal_114;

  reg [2:0] rvx_signal_172;

  reg [2:0] rvx_signal_266;

  reg [2:0] rvx_signal_444;

  reg [2:0] rvx_signal_088;

  reg [2:0] rvx_signal_234;

  reg [2:0] rvx_signal_097;

  reg [2:0] rvx_signal_267;

  reg [2:0] rvx_signal_248;

  reg [2:0] rvx_signal_400;

  reg [2:0] rvx_signal_430;

  reg [2:0] rvx_signal_359;

  reg [2:0] rvx_signal_332;

  reg [2:0] rvx_signal_300;

  reg [2:0] rvx_signal_032;

  reg [2:0] rvx_signal_435;

  reg  rvx_signal_065;

  reg  rvx_signal_437;

  reg  rvx_signal_382;

  reg  rvx_signal_316;

  reg  rvx_signal_165;

  reg  rvx_signal_004;

  reg  rvx_signal_272;

  reg  rvx_signal_409;

  reg  rvx_signal_202;

  reg  rvx_signal_454;

  reg  rvx_signal_092;

  reg  rvx_signal_298;

  reg  rvx_signal_096;

  reg  rvx_signal_167;

  reg  rvx_signal_294;

  reg  rvx_signal_371;

  reg  rvx_signal_103;

  reg  rvx_signal_019;

  reg  rvx_signal_080;

  reg  rvx_signal_239;

  reg  rvx_signal_124;

  reg  rvx_signal_222;

  reg  rvx_signal_306;

  reg  rvx_signal_238;

  reg  rvx_signal_011;

  reg  rvx_signal_029;

  reg  rvx_signal_166;

  reg  rvx_signal_228;

  reg  rvx_signal_183;

  reg  rvx_signal_253;

  reg  rvx_signal_033;

  reg  rvx_signal_229;

  reg  rvx_signal_099;

  reg  rvx_signal_369;

  reg  rvx_signal_221;

  reg  rvx_signal_224;

  reg  rvx_signal_066;

  reg  rvx_signal_111;

  reg  rvx_signal_179;

  reg  rvx_signal_050;

  reg  rvx_signal_215;

  reg  rvx_signal_386;

  reg  rvx_signal_450;

  reg  rvx_signal_399;

  reg  rvx_signal_067;

  reg  rvx_signal_350;

  reg  rvx_signal_265;

  reg  rvx_signal_304;

  reg  rvx_signal_058;

  reg  rvx_signal_433;

  reg  rvx_signal_465;

  reg  rvx_signal_197;

  reg  rvx_signal_358;

  reg  rvx_signal_436;

  reg  rvx_signal_001;

  reg  rvx_signal_131;

  reg  rvx_signal_410;

  reg  rvx_signal_137;

  reg  rvx_signal_178;

  reg  rvx_signal_052;

  reg  rvx_signal_423;

  reg  rvx_signal_462;

  reg  rvx_signal_475;

  reg  rvx_signal_408;

  reg [5:0] rvx_signal_153;

  wire  _T_1259;
  wire [3:0] _T_1260;
  wire  _T_1261;
  wire [3:0] _T_1262;
  wire  _T_1263;
  wire [3:0] _T_1264;
  wire  _T_1265;
  wire [3:0] _T_1266;
  wire  _T_1267;
  wire [3:0] _T_1268;
  wire  _T_1269;
  wire [3:0] _T_1270;
  wire  _T_1271;
  wire [3:0] _T_1272;
  wire  _T_1273;
  wire [3:0] _T_1274;
  wire  _T_1275;
  wire [3:0] _T_1276;
  wire  _T_1277;
  wire [3:0] _T_1278;
  wire  _T_1279;
  wire [3:0] _T_1280;
  wire  _T_1281;
  wire [3:0] _T_1282;
  wire  _T_1283;
  wire [3:0] _T_1284;
  wire  _T_1285;
  wire [3:0] _T_1286;
  wire  _T_1287;
  wire [3:0] _T_1288;
  wire  _T_1289;
  wire [3:0] _T_1290;
  wire  _T_1291;
  wire [3:0] _T_1292;
  wire  _T_1293;
  wire [3:0] _T_1294;
  wire  _T_1295;
  wire [3:0] _T_1296;
  wire  _T_1297;
  wire [3:0] _T_1298;
  wire  _T_1299;
  wire [3:0] _T_1300;
  wire  _T_1301;
  wire [3:0] _T_1302;
  wire  _T_1303;
  wire [3:0] _T_1304;
  wire  _T_1305;
  wire [3:0] _T_1306;
  wire  _T_1307;
  wire [3:0] _T_1308;
  wire  _T_1309;
  wire [3:0] _T_1310;
  wire  _T_1311;
  wire [3:0] _T_1312;
  wire  _T_1313;
  wire [3:0] _T_1314;
  wire  _T_1315;
  wire [3:0] _T_1316;
  wire  _T_1317;
  wire [3:0] _T_1318;
  wire  _T_1319;
  wire [3:0] _T_1320;
  wire  _T_1321;
  wire [3:0] _T_1322;
  wire  _T_1325;
  wire [3:0] _T_1328;
  wire  _T_1329;
  wire  _T_1332;
  wire [3:0] _T_1335;
  wire  _T_1336;
  wire  _T_1337;
  wire [1:0] _GEN_3205;
  wire [1:0] _T_1339;
  wire [3:0] _T_1340;
  wire [1:0] _T_1341;
  wire  _T_1344;
  wire [3:0] _T_1347;
  wire  _T_1348;
  wire  _T_1351;
  wire [3:0] _T_1354;
  wire  _T_1355;
  wire  _T_1356;
  wire [1:0] _GEN_3206;
  wire [1:0] _T_1358;
  wire [3:0] _T_1359;
  wire [1:0] _T_1360;
  wire  _T_1361;
  wire [2:0] _GEN_3207;
  wire [2:0] _T_1363;
  wire [3:0] _T_1364;
  wire [2:0] _T_1365;
  wire  _T_1368;
  wire [3:0] _T_1371;
  wire  _T_1372;
  wire  _T_1375;
  wire [3:0] _T_1378;
  wire  _T_1379;
  wire  _T_1380;
  wire [1:0] _GEN_3208;
  wire [1:0] _T_1382;
  wire [3:0] _T_1383;
  wire [1:0] _T_1384;
  wire  _T_1387;
  wire [3:0] _T_1390;
  wire  _T_1391;
  wire  _T_1394;
  wire [3:0] _T_1397;
  wire  _T_1398;
  wire  _T_1399;
  wire [1:0] _GEN_3209;
  wire [1:0] _T_1401;
  wire [3:0] _T_1402;
  wire [1:0] _T_1403;
  wire  _T_1404;
  wire [2:0] _GEN_3210;
  wire [2:0] _T_1406;
  wire [3:0] _T_1407;
  wire [2:0] _T_1408;
  wire  _T_1409;
  wire [3:0] _GEN_3211;
  wire [3:0] _T_1411;
  wire [3:0] _T_1412;
  wire [3:0] _T_1413;
  wire  _T_1416;
  wire [3:0] _T_1419;
  wire  _T_1420;
  wire  _T_1423;
  wire [3:0] _T_1426;
  wire  _T_1427;
  wire  _T_1428;
  wire [1:0] _GEN_3212;
  wire [1:0] _T_1430;
  wire [3:0] _T_1431;
  wire [1:0] _T_1432;
  wire  _T_1435;
  wire [3:0] _T_1438;
  wire  _T_1439;
  wire  _T_1442;
  wire [3:0] _T_1445;
  wire  _T_1446;
  wire  _T_1447;
  wire [1:0] _GEN_3213;
  wire [1:0] _T_1449;
  wire [3:0] _T_1450;
  wire [1:0] _T_1451;
  wire  _T_1452;
  wire [2:0] _GEN_3214;
  wire [2:0] _T_1454;
  wire [3:0] _T_1455;
  wire [2:0] _T_1456;
  wire  _T_1459;
  wire [3:0] _T_1462;
  wire  _T_1463;
  wire  _T_1466;
  wire [3:0] _T_1469;
  wire  _T_1470;
  wire  _T_1471;
  wire [1:0] _GEN_3215;
  wire [1:0] _T_1473;
  wire [3:0] _T_1474;
  wire [1:0] _T_1475;
  wire  _T_1478;
  wire [3:0] _T_1481;
  wire  _T_1482;
  wire  _T_1485;
  wire [3:0] _T_1488;
  wire  _T_1489;
  wire  _T_1490;
  wire [1:0] _GEN_3216;
  wire [1:0] _T_1492;
  wire [3:0] _T_1493;
  wire [1:0] _T_1494;
  wire  _T_1495;
  wire [2:0] _GEN_3217;
  wire [2:0] _T_1497;
  wire [3:0] _T_1498;
  wire [2:0] _T_1499;
  wire  _T_1500;
  wire [3:0] _GEN_3218;
  wire [3:0] _T_1502;
  wire [3:0] _T_1503;
  wire [3:0] _T_1504;
  wire  _T_1505;
  wire [4:0] _GEN_3219;
  wire [4:0] _T_1507;
  wire [3:0] _T_1508;
  wire [4:0] _T_1509;
  wire  _T_1511;
  wire [3:0] _T_1514;
  wire [5:0] _T_1515;
  reg [3:0] _T_1517;

  wire [3:0] _T_1519;
  wire  _T_1520;
  wire  rvx_signal_189;
  wire [1:0] _T_1529;
  wire [1:0] _T_1530;
  wire  _T_1531;
  wire  _T_1532;
  wire  _T_1534;
  wire  _T_1536;
  wire  _T_1538;
  wire [63:0] _T_1541;
  wire [32:0] _T_1542;
  wire [32:0] _T_1544;
  wire [32:0] rvx_signal_161;
  wire  _T_1551;
  wire  _T_1552;
  wire  _T_1553;
  wire  _T_1554;
  wire  _T_1555;
  wire  _T_1556;
  wire  _T_1557;
  wire  _T_1558;
  wire  _T_1559;
  wire  _T_1560;
  wire  _T_1561;
  wire  _T_1562;
  wire  _T_1563;
  wire  _T_1564;
  wire  _T_1565;
  wire  _T_1566;
  wire  _T_1567;
  wire  _T_1568;
  wire  _T_1569;
  wire  _T_1570;
  wire  _T_1571;
  wire  _T_1572;
  wire  _T_1573;
  wire  _T_1574;
  wire  _T_1575;
  wire  _T_1576;
  wire  _T_1577;
  wire  _T_1578;
  wire  _T_1579;
  wire  _T_1580;
  wire  _T_1581;
  wire  _T_1582;
  wire  rvx_signal_017;
  wire  rvx_signal_164;
  wire  rvx_signal_427;
  wire  rvx_signal_005;
  wire  rvx_signal_275;
  wire  rvx_signal_182;
  wire  rvx_signal_185;
  wire  rvx_signal_110;
  wire  rvx_signal_372;
  wire  rvx_signal_290;
  wire  rvx_signal_407;
  wire  rvx_signal_126;
  wire  rvx_signal_374;
  wire  rvx_signal_318;
  wire  rvx_signal_279;
  wire  rvx_signal_303;
  wire  rvx_signal_038;
  wire  rvx_signal_077;
  wire  rvx_signal_384;
  wire  rvx_signal_446;
  wire  rvx_signal_443;
  wire  rvx_signal_150;
  wire  rvx_signal_383;
  wire  rvx_signal_048;
  wire  rvx_signal_249;
  wire  rvx_signal_064;
  wire  rvx_signal_470;
  wire  rvx_signal_258;
  wire  rvx_signal_034;
  wire  rvx_signal_018;
  wire  rvx_signal_155;
  wire  rvx_signal_144;
  wire  _T_1626;
  wire  _T_1627;
  wire  _T_1629;
  wire  _GEN_8;
  wire  _T_1631;
  wire  _T_1632;
  wire  _T_1634;
  wire  _GEN_9;
  wire  _T_1636;
  wire  _T_1637;
  wire  _T_1639;
  wire  _GEN_10;
  wire  _T_1641;
  wire  _T_1642;
  wire  _T_1644;
  wire  _GEN_11;
  wire  _T_1646;
  wire  _T_1647;
  wire  _T_1649;
  wire  _GEN_12;
  wire  _T_1651;
  wire  _T_1652;
  wire  _T_1654;
  wire  _GEN_13;
  wire  _T_1656;
  wire  _T_1657;
  wire  _T_1659;
  wire  _GEN_14;
  wire  _T_1661;
  wire  _T_1662;
  wire  _T_1664;
  wire  _GEN_15;
  wire  _T_1666;
  wire  _T_1667;
  wire  _T_1669;
  wire  _GEN_16;
  wire  _T_1671;
  wire  _T_1672;
  wire  _T_1674;
  wire  _GEN_17;
  wire  _T_1676;
  wire  _T_1677;
  wire  _T_1679;
  wire  _GEN_18;
  wire  _T_1681;
  wire  _T_1682;
  wire  _T_1684;
  wire  _GEN_19;
  wire  _T_1686;
  wire  _T_1687;
  wire  _T_1689;
  wire  _GEN_20;
  wire  _T_1691;
  wire  _T_1692;
  wire  _T_1694;
  wire  _GEN_21;
  wire  _T_1696;
  wire  _T_1697;
  wire  _T_1699;
  wire  _GEN_22;
  wire  _T_1701;
  wire  _T_1702;
  wire  _T_1704;
  wire  _GEN_23;
  wire  _T_1706;
  wire  _T_1707;
  wire  _T_1709;
  wire  _GEN_24;
  wire  _T_1711;
  wire  _T_1712;
  wire  _T_1714;
  wire  _GEN_25;
  wire  _T_1716;
  wire  _T_1717;
  wire  _T_1719;
  wire  _GEN_26;
  wire  _T_1721;
  wire  _T_1722;
  wire  _T_1724;
  wire  _GEN_27;
  wire  _T_1726;
  wire  _T_1727;
  wire  _T_1729;
  wire  _GEN_28;
  wire  _T_1731;
  wire  _T_1732;
  wire  _T_1734;
  wire  _GEN_29;
  wire  _T_1736;
  wire  _T_1737;
  wire  _T_1739;
  wire  _GEN_30;
  wire  _T_1741;
  wire  _T_1742;
  wire  _T_1744;
  wire  _GEN_31;
  wire  _T_1746;
  wire  _T_1747;
  wire  _T_1749;
  wire  _GEN_32;
  wire  _T_1751;
  wire  _T_1752;
  wire  _T_1754;
  wire  _GEN_33;
  wire  _T_1756;
  wire  _T_1757;
  wire  _T_1759;
  wire  _GEN_34;
  wire  _T_1761;
  wire  _T_1762;
  wire  _T_1764;
  wire  _GEN_35;
  wire  _T_1766;
  wire  _T_1767;
  wire  _T_1769;
  wire  _GEN_36;
  wire  _T_1771;
  wire  _T_1772;
  wire  _T_1774;
  wire  _GEN_37;
  wire  _T_1776;
  wire  _T_1777;
  wire  _T_1779;
  wire  _GEN_38;
  wire  _T_1781;
  wire  _T_1782;
  wire  _T_1784;
  wire  _GEN_39;
  wire  rvx_signal_431;
  wire [1:0] _T_1792;
  wire [1:0] _T_1793;
  wire  _T_1794;
  wire  _T_1795;
  wire  _T_1797;
  wire  _T_1799;
  wire  _T_1801;
  wire [5:0] rvx_signal_120;
  wire [63:0] _T_1805;
  wire [32:0] _T_1806;
  wire [32:0] rvx_signal_432;
  wire  _T_1808;
  wire  _T_1809;
  wire  _T_1810;
  wire  _T_1811;
  wire  _T_1812;
  wire  _T_1813;
  wire  _T_1814;
  wire  _T_1815;
  wire  _T_1816;
  wire  _T_1817;
  wire  _T_1818;
  wire  _T_1819;
  wire  _T_1820;
  wire  _T_1821;
  wire  _T_1822;
  wire  _T_1823;
  wire  _T_1824;
  wire  _T_1825;
  wire  _T_1826;
  wire  _T_1827;
  wire  _T_1828;
  wire  _T_1829;
  wire  _T_1830;
  wire  _T_1831;
  wire  _T_1832;
  wire  _T_1833;
  wire  _T_1834;
  wire  _T_1835;
  wire  _T_1836;
  wire  _T_1837;
  wire  _T_1838;
  wire  _T_1839;
  wire  _T_1840;
  wire  _T_1846_ready;
  wire  _T_1846_valid;
  wire  _T_1846_bits_read;
  wire [23:0] _T_1846_bits_index;
  wire [31:0] _T_1846_bits_data;
  wire [3:0] _T_1846_bits_mask;
  wire [11:0] _T_1846_bits_extra;
  wire  _T_1851;
  wire [25:0] _T_1852;
  wire [11:0] _T_1853;
  wire  _T_1859_ready;
  wire  _T_1859_valid;
  wire  _T_1859_bits_read;
  wire [31:0] _T_1859_bits_data;
  wire [11:0] _T_1859_bits_extra;
  wire  _T_1868_ready;
  wire  _T_1868_valid;
  wire  _T_1868_bits_read;
  wire [23:0] _T_1868_bits_index;
  wire [31:0] _T_1868_bits_data;
  wire [3:0] _T_1868_bits_mask;
  wire [11:0] _T_1868_bits_extra;
  wire  rvx_signal_043;
  wire  rvx_signal_242;
  wire  rvx_signal_296;
  wire  rvx_signal_007;
  wire  rvx_signal_255;
  wire [23:0] rvx_signal_364;
  wire [31:0] rvx_signal_129;
  wire [3:0] rvx_signal_045;
  wire [11:0] rvx_signal_240;
  wire  rvx_signal_426;
  wire  rvx_signal_309;
  wire  rvx_signal_388;
  wire [23:0] rvx_signal_060;
  wire [31:0] rvx_signal_162;
  wire [3:0] rvx_signal_429;
  wire [11:0] rvx_signal_263;
  wire [23:0] _T_2903;
  wire [23:0] _T_2904;
  wire  _T_2906;
  wire [23:0] _T_2912;
  wire [23:0] _T_2913;
  wire  _T_2915;
  wire [23:0] _T_2921;
  wire [23:0] _T_2922;
  wire  _T_2924;
  wire [23:0] _T_2930;
  wire [23:0] _T_2931;
  wire  _T_2933;
  wire [23:0] _T_2939;
  wire [23:0] _T_2940;
  wire  _T_2942;
  wire [23:0] _T_2948;
  wire [23:0] _T_2949;
  wire  _T_2951;
  wire [23:0] _T_2957;
  wire [23:0] _T_2958;
  wire  _T_2960;
  wire [23:0] _T_2966;
  wire [23:0] _T_2967;
  wire  _T_2969;
  wire [23:0] _T_2975;
  wire [23:0] _T_2976;
  wire  _T_2978;
  wire [23:0] _T_2984;
  wire [23:0] _T_2985;
  wire  _T_2987;
  wire [23:0] _T_2993;
  wire [23:0] _T_2994;
  wire  _T_2996;
  wire [23:0] _T_3002;
  wire [23:0] _T_3003;
  wire  _T_3005;
  wire [23:0] _T_3011;
  wire [23:0] _T_3012;
  wire  _T_3014;
  wire [23:0] _T_3020;
  wire [23:0] _T_3021;
  wire  _T_3023;
  wire [23:0] _T_3029;
  wire [23:0] _T_3030;
  wire  _T_3032;
  wire [23:0] _T_3038;
  wire [23:0] _T_3039;
  wire  _T_3041;
  wire [23:0] _T_3047;
  wire [23:0] _T_3048;
  wire  _T_3050;
  wire [23:0] _T_3056;
  wire [23:0] _T_3057;
  wire  _T_3059;
  wire [23:0] _T_3065;
  wire [23:0] _T_3066;
  wire  _T_3068;
  wire [23:0] _T_3074;
  wire [23:0] _T_3075;
  wire  _T_3077;
  wire [23:0] _T_3083;
  wire [23:0] _T_3084;
  wire  _T_3086;
  wire [23:0] _T_3092;
  wire [23:0] _T_3093;
  wire  _T_3095;
  wire [23:0] _T_3101;
  wire [23:0] _T_3102;
  wire  _T_3104;
  wire [23:0] _T_3110;
  wire [23:0] _T_3111;
  wire  _T_3113;
  wire [23:0] _T_3119;
  wire [23:0] _T_3120;
  wire  _T_3122;
  wire [23:0] _T_3128;
  wire [23:0] _T_3129;
  wire  _T_3131;
  wire [23:0] _T_3137;
  wire [23:0] _T_3138;
  wire  _T_3140;
  wire [23:0] _T_3146;
  wire [23:0] _T_3147;
  wire  _T_3149;
  wire [23:0] _T_3155;
  wire [23:0] _T_3156;
  wire  _T_3158;
  wire [23:0] _T_3164;
  wire [23:0] _T_3165;
  wire  _T_3167;
  wire [23:0] _T_3173;
  wire [23:0] _T_3174;
  wire  _T_3176;
  wire [23:0] _T_3182;
  wire [23:0] _T_3183;
  wire  _T_3185;
  wire [23:0] _T_3191;
  wire [23:0] _T_3192;
  wire  _T_3194;
  wire [23:0] _T_3200;
  wire [23:0] _T_3201;
  wire  _T_3203;
  wire [23:0] _T_3209;
  wire [23:0] _T_3210;
  wire  _T_3212;
  wire [23:0] _T_3218;
  wire [23:0] _T_3219;
  wire  _T_3221;
  wire [23:0] _T_3227;
  wire [23:0] _T_3228;
  wire  _T_3230;
  wire [23:0] _T_3236;
  wire [23:0] _T_3237;
  wire  _T_3239;
  wire [23:0] _T_3245;
  wire [23:0] _T_3246;
  wire  _T_3248;
  wire  _T_3466_41;
  wire  _T_3573_33;
  wire  _T_3573_34;
  wire  _T_3573_35;
  wire  _T_3573_36;
  wire  _T_3573_37;
  wire  _T_3573_38;
  wire  _T_3573_39;
  wire  _T_3573_40;
  wire  _T_3573_41;
  wire  _T_3573_42;
  wire  _T_3573_43;
  wire  _T_3573_44;
  wire  _T_3573_45;
  wire  _T_3573_46;
  wire  _T_3573_47;
  wire  _T_3573_48;
  wire  _T_3573_49;
  wire  _T_3573_50;
  wire  _T_3573_51;
  wire  _T_3573_53;
  wire  _T_3573_54;
  wire  _T_3573_55;
  wire  _T_3573_56;
  wire  _T_3573_57;
  wire  _T_3573_58;
  wire  _T_3573_59;
  wire  _T_3573_60;
  wire  _T_3573_61;
  wire  _T_3573_62;
  wire  _T_3573_63;
  wire  _T_3573_64;
  wire  _T_3573_65;
  wire  _T_3573_66;
  wire  _T_3573_67;
  wire  _T_3573_68;
  wire  _T_3573_69;
  wire  _T_3573_70;
  wire  _T_3573_71;
  wire  _T_3573_72;
  wire  _T_3573_73;
  wire  _T_3573_74;
  wire  _T_3573_75;
  wire  _T_3573_76;
  wire  _T_3573_77;
  wire  _T_3573_78;
  wire  _T_3573_79;
  wire  _T_3573_80;
  wire  _T_3573_81;
  wire  _T_3573_82;
  wire  _T_3573_83;
  wire  _T_3573_84;
  wire  _T_3573_85;
  wire  _T_3573_86;
  wire  _T_3573_87;
  wire  _T_3573_88;
  wire  _T_3573_90;
  wire  _T_3573_91;
  wire  _T_3573_92;
  wire  _T_3573_93;
  wire  _T_3573_94;
  wire  _T_3573_95;
  wire  _T_3573_96;
  wire  _T_3573_97;
  wire  _T_3573_98;
  wire  _T_3573_99;
  wire  _T_3573_100;
  wire  _T_4212;
  wire  _T_4213;
  wire  _T_4214;
  wire  _T_4215;
  wire [7:0] _T_4219;
  wire [7:0] _T_4223;
  wire [7:0] _T_4227;
  wire [7:0] _T_4231;
  wire [15:0] _T_4232;
  wire [15:0] _T_4233;
  wire [31:0] _T_4234;
  wire  _T_4242;
  wire  _T_4246;
  wire  _T_4248;
  wire  _T_4255;
  wire  _T_4282;
  wire  _T_4286;
  wire  _T_4288;
  wire  _T_4295;
  wire [1:0] _GEN_3220;
  wire [1:0] _T_4310;
  wire  _T_4322;
  wire  _T_4326;
  wire  _T_4328;
  wire  _T_4335;
  wire [2:0] _GEN_3221;
  wire [2:0] _T_4350;
  wire [2:0] _GEN_3222;
  wire [2:0] _T_4354;
  wire  _T_4362;
  wire  _T_4366;
  wire  _T_4368;
  wire  _T_4375;
  wire [3:0] _GEN_3223;
  wire [3:0] _T_4390;
  wire [3:0] _GEN_3224;
  wire [3:0] _T_4394;
  wire  _T_4402;
  wire  _T_4406;
  wire  _T_4408;
  wire  _T_4415;
  wire [4:0] _GEN_3225;
  wire [4:0] _T_4430;
  wire [4:0] _GEN_3226;
  wire [4:0] _T_4434;
  wire  _T_4442;
  wire  _T_4446;
  wire  _T_4448;
  wire  _T_4455;
  wire [5:0] _GEN_3227;
  wire [5:0] _T_4470;
  wire [5:0] _GEN_3228;
  wire [5:0] _T_4474;
  wire  _T_4482;
  wire  _T_4486;
  wire  _T_4488;
  wire  _T_4495;
  wire [6:0] _GEN_3229;
  wire [6:0] _T_4510;
  wire [6:0] _GEN_3230;
  wire [6:0] _T_4514;
  wire  _T_4522;
  wire  _T_4526;
  wire  _T_4528;
  wire  _T_4535;
  wire [7:0] _GEN_3231;
  wire [7:0] _T_4550;
  wire [7:0] _GEN_3232;
  wire [7:0] _T_4554;
  wire  _T_4562;
  wire  _T_4566;
  wire  _T_4568;
  wire  _T_4575;
  wire [8:0] _GEN_3233;
  wire [8:0] _T_4590;
  wire [8:0] _GEN_3234;
  wire [8:0] _T_4594;
  wire  _T_4602;
  wire  _T_4606;
  wire  _T_4608;
  wire  _T_4615;
  wire [9:0] _GEN_3235;
  wire [9:0] _T_4630;
  wire [9:0] _GEN_3236;
  wire [9:0] _T_4634;
  wire  _T_4642;
  wire  _T_4646;
  wire  _T_4648;
  wire  _T_4655;
  wire [10:0] _GEN_3237;
  wire [10:0] _T_4670;
  wire [10:0] _GEN_3238;
  wire [10:0] _T_4674;
  wire  _T_4682;
  wire  _T_4686;
  wire  _T_4688;
  wire  _T_4695;
  wire [11:0] _GEN_3239;
  wire [11:0] _T_4710;
  wire [11:0] _GEN_3240;
  wire [11:0] _T_4714;
  wire  _T_4722;
  wire  _T_4726;
  wire  _T_4728;
  wire  _T_4735;
  wire [12:0] _GEN_3241;
  wire [12:0] _T_4750;
  wire [12:0] _GEN_3242;
  wire [12:0] _T_4754;
  wire  _T_4762;
  wire  _T_4766;
  wire  _T_4768;
  wire  _T_4775;
  wire [13:0] _GEN_3243;
  wire [13:0] _T_4790;
  wire [13:0] _GEN_3244;
  wire [13:0] _T_4794;
  wire  _T_4802;
  wire  _T_4806;
  wire  _T_4808;
  wire  _T_4815;
  wire [14:0] _GEN_3245;
  wire [14:0] _T_4830;
  wire [14:0] _GEN_3246;
  wire [14:0] _T_4834;
  wire  _T_4842;
  wire  _T_4846;
  wire  _T_4848;
  wire  _T_4855;
  wire [15:0] _GEN_3247;
  wire [15:0] _T_4870;
  wire [15:0] _GEN_3248;
  wire [15:0] _T_4874;
  wire  _T_4882;
  wire  _T_4886;
  wire  _T_4888;
  wire  _T_4895;
  wire [16:0] _GEN_3249;
  wire [16:0] _T_4910;
  wire [16:0] _GEN_3250;
  wire [16:0] _T_4914;
  wire  _T_4922;
  wire  _T_4926;
  wire  _T_4928;
  wire  _T_4935;
  wire [17:0] _GEN_3251;
  wire [17:0] _T_4950;
  wire [17:0] _GEN_3252;
  wire [17:0] _T_4954;
  wire  _T_4962;
  wire  _T_4966;
  wire  _T_4968;
  wire  _T_4975;
  wire [18:0] _GEN_3253;
  wire [18:0] _T_4990;
  wire [18:0] _GEN_3254;
  wire [18:0] _T_4994;
  wire  _T_5002;
  wire  _T_5006;
  wire  _T_5008;
  wire  _T_5015;
  wire [19:0] _GEN_3255;
  wire [19:0] _T_5030;
  wire [19:0] _GEN_3256;
  wire [19:0] _T_5034;
  wire  _T_5042;
  wire  _T_5046;
  wire  _T_5048;
  wire  _T_5055;
  wire [20:0] _GEN_3257;
  wire [20:0] _T_5070;
  wire [20:0] _GEN_3258;
  wire [20:0] _T_5074;
  wire  _T_5082;
  wire  _T_5086;
  wire  _T_5088;
  wire  _T_5095;
  wire [21:0] _GEN_3259;
  wire [21:0] _T_5110;
  wire [21:0] _GEN_3260;
  wire [21:0] _T_5114;
  wire  _T_5122;
  wire  _T_5126;
  wire  _T_5128;
  wire  _T_5135;
  wire [22:0] _GEN_3261;
  wire [22:0] _T_5150;
  wire [22:0] _GEN_3262;
  wire [22:0] _T_5154;
  wire  _T_5162;
  wire  _T_5166;
  wire  _T_5168;
  wire  _T_5175;
  wire [23:0] _GEN_3263;
  wire [23:0] _T_5190;
  wire [23:0] _GEN_3264;
  wire [23:0] _T_5194;
  wire  _T_5202;
  wire  _T_5206;
  wire  _T_5208;
  wire  _T_5215;
  wire [24:0] _GEN_3265;
  wire [24:0] _T_5230;
  wire [24:0] _GEN_3266;
  wire [24:0] _T_5234;
  wire  _T_5242;
  wire  _T_5246;
  wire  _T_5248;
  wire  _T_5255;
  wire [25:0] _GEN_3267;
  wire [25:0] _T_5270;
  wire [25:0] _GEN_3268;
  wire [25:0] _T_5274;
  wire  _T_5282;
  wire  _T_5286;
  wire  _T_5288;
  wire  _T_5295;
  wire [26:0] _GEN_3269;
  wire [26:0] _T_5310;
  wire [26:0] _GEN_3270;
  wire [26:0] _T_5314;
  wire  _T_5322;
  wire  _T_5326;
  wire  _T_5328;
  wire  _T_5335;
  wire [27:0] _GEN_3271;
  wire [27:0] _T_5350;
  wire [27:0] _GEN_3272;
  wire [27:0] _T_5354;
  wire  _T_5362;
  wire  _T_5366;
  wire  _T_5368;
  wire  _T_5375;
  wire [28:0] _GEN_3273;
  wire [28:0] _T_5390;
  wire [28:0] _GEN_3274;
  wire [28:0] _T_5394;
  wire  _T_5402;
  wire  _T_5406;
  wire  _T_5408;
  wire  _T_5415;
  wire [29:0] _GEN_3275;
  wire [29:0] _T_5430;
  wire [29:0] _GEN_3276;
  wire [29:0] _T_5434;
  wire  _T_5442;
  wire  _T_5446;
  wire  _T_5448;
  wire  _T_5455;
  wire [30:0] _GEN_3277;
  wire [30:0] _T_5470;
  wire [30:0] _GEN_3278;
  wire [30:0] _T_5474;
  wire  _T_5482;
  wire  _T_5486;
  wire  _T_5488;
  wire  _T_5495;
  wire [31:0] _GEN_3279;
  wire [31:0] _T_5510;
  wire [31:0] _GEN_3280;
  wire [31:0] _T_5514;
  wire  _T_5524;
  wire [31:0] _T_5526;
  wire  _T_5528;
  wire [31:0] _T_5535;
  wire  _T_5574;
  wire [31:0] _GEN_41;
  wire [31:0] _T_5593;
  wire  _T_5614;
  wire [31:0] _GEN_42;
  wire [31:0] _T_5633;
  wire  _T_5654;
  wire [31:0] _GEN_43;
  wire [31:0] _T_5673;
  wire  _T_5694;
  wire [31:0] _GEN_44;
  wire [31:0] _T_5713;
  wire  _T_5734;
  wire [31:0] _GEN_45;
  wire [31:0] _T_5753;
  wire  _T_5774;
  wire [31:0] _GEN_46;
  wire [31:0] _T_5793;
  wire  _T_5814;
  wire  _GEN_47;
  wire  _T_5854;
  wire [31:0] _GEN_48;
  wire [31:0] _T_5873;
  wire  _T_5890;
  wire  _T_5894;
  wire [5:0] _T_5897;
  wire  _T_5898;
  wire  _T_5900;
  wire  _T_5902;
  wire  _GEN_0;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _T_5906;
  wire [31:0] _T_5923;
  wire  _T_5944;
  wire [31:0] _GEN_81;
  wire [31:0] _T_5963;
  wire  _T_5984;
  wire [31:0] _GEN_82;
  wire [31:0] _T_6003;
  wire  _T_6024;
  wire [31:0] _GEN_83;
  wire [31:0] _T_6043;
  wire  _T_6064;
  wire [31:0] _GEN_84;
  wire [31:0] _T_6083;
  wire  _T_6104;
  wire [31:0] _GEN_85;
  wire [31:0] _T_6123;
  wire  _T_6144;
  wire [31:0] _GEN_86;
  wire [31:0] _T_6163;
  wire  _T_6184;
  wire [31:0] _GEN_87;
  wire [31:0] _T_6203;
  wire  _T_6224;
  wire [31:0] _GEN_88;
  wire [31:0] _T_6243;
  wire  _T_6264;
  wire [31:0] _GEN_89;
  wire [31:0] _T_6283;
  wire  _T_6304;
  wire [31:0] _GEN_90;
  wire [31:0] _T_6323;
  wire  _T_6384;
  wire  _GEN_92;
  wire [1:0] _GEN_3281;
  wire [1:0] _T_6400;
  wire  _T_6424;
  wire  _GEN_93;
  wire [2:0] _GEN_3282;
  wire [2:0] _T_6440;
  wire [2:0] _GEN_3283;
  wire [2:0] _T_6444;
  wire  _T_6464;
  wire  _GEN_94;
  wire [3:0] _GEN_3284;
  wire [3:0] _T_6480;
  wire [3:0] _GEN_3285;
  wire [3:0] _T_6484;
  wire  _T_6504;
  wire  _GEN_95;
  wire [4:0] _GEN_3286;
  wire [4:0] _T_6520;
  wire [4:0] _GEN_3287;
  wire [4:0] _T_6524;
  wire  _T_6544;
  wire  _GEN_96;
  wire [5:0] _GEN_3288;
  wire [5:0] _T_6560;
  wire [5:0] _GEN_3289;
  wire [5:0] _T_6564;
  wire  _T_6584;
  wire  _GEN_97;
  wire [6:0] _GEN_3290;
  wire [6:0] _T_6600;
  wire [6:0] _GEN_3291;
  wire [6:0] _T_6604;
  wire  _T_6624;
  wire  _GEN_98;
  wire [7:0] _GEN_3292;
  wire [7:0] _T_6640;
  wire [7:0] _GEN_3293;
  wire [7:0] _T_6644;
  wire  _T_6664;
  wire  _GEN_99;
  wire [8:0] _GEN_3294;
  wire [8:0] _T_6680;
  wire [8:0] _GEN_3295;
  wire [8:0] _T_6684;
  wire  _T_6704;
  wire  _GEN_100;
  wire [9:0] _GEN_3296;
  wire [9:0] _T_6720;
  wire [9:0] _GEN_3297;
  wire [9:0] _T_6724;
  wire  _T_6744;
  wire  _GEN_101;
  wire [10:0] _GEN_3298;
  wire [10:0] _T_6760;
  wire [10:0] _GEN_3299;
  wire [10:0] _T_6764;
  wire  _T_6784;
  wire  _GEN_102;
  wire [11:0] _GEN_3300;
  wire [11:0] _T_6800;
  wire [11:0] _GEN_3301;
  wire [11:0] _T_6804;
  wire  _T_6824;
  wire  _GEN_103;
  wire [12:0] _GEN_3302;
  wire [12:0] _T_6840;
  wire [12:0] _GEN_3303;
  wire [12:0] _T_6844;
  wire  _T_6864;
  wire  _GEN_104;
  wire [13:0] _GEN_3304;
  wire [13:0] _T_6880;
  wire [13:0] _GEN_3305;
  wire [13:0] _T_6884;
  wire  _T_6904;
  wire  _GEN_105;
  wire [14:0] _GEN_3306;
  wire [14:0] _T_6920;
  wire [14:0] _GEN_3307;
  wire [14:0] _T_6924;
  wire  _T_6944;
  wire  _GEN_106;
  wire [15:0] _GEN_3308;
  wire [15:0] _T_6960;
  wire [15:0] _GEN_3309;
  wire [15:0] _T_6964;
  wire  _T_6984;
  wire  _GEN_107;
  wire [16:0] _GEN_3310;
  wire [16:0] _T_7000;
  wire [16:0] _GEN_3311;
  wire [16:0] _T_7004;
  wire  _T_7024;
  wire  _GEN_108;
  wire [17:0] _GEN_3312;
  wire [17:0] _T_7040;
  wire [17:0] _GEN_3313;
  wire [17:0] _T_7044;
  wire  _T_7064;
  wire  _GEN_109;
  wire [18:0] _GEN_3314;
  wire [18:0] _T_7080;
  wire [18:0] _GEN_3315;
  wire [18:0] _T_7084;
  wire  _T_7104;
  wire  _GEN_110;
  wire [19:0] _GEN_3316;
  wire [19:0] _T_7120;
  wire [19:0] _GEN_3317;
  wire [19:0] _T_7124;
  wire  _T_7144;
  wire  _GEN_111;
  wire [20:0] _GEN_3318;
  wire [20:0] _T_7160;
  wire [20:0] _GEN_3319;
  wire [20:0] _T_7164;
  wire  _T_7184;
  wire  _GEN_112;
  wire [21:0] _GEN_3320;
  wire [21:0] _T_7200;
  wire [21:0] _GEN_3321;
  wire [21:0] _T_7204;
  wire  _T_7224;
  wire  _GEN_113;
  wire [22:0] _GEN_3322;
  wire [22:0] _T_7240;
  wire [22:0] _GEN_3323;
  wire [22:0] _T_7244;
  wire  _T_7264;
  wire  _GEN_114;
  wire [23:0] _GEN_3324;
  wire [23:0] _T_7280;
  wire [23:0] _GEN_3325;
  wire [23:0] _T_7284;
  wire  _T_7304;
  wire  _GEN_115;
  wire [24:0] _GEN_3326;
  wire [24:0] _T_7320;
  wire [24:0] _GEN_3327;
  wire [24:0] _T_7324;
  wire  _T_7344;
  wire  _GEN_116;
  wire [25:0] _GEN_3328;
  wire [25:0] _T_7360;
  wire [25:0] _GEN_3329;
  wire [25:0] _T_7364;
  wire  _T_7384;
  wire  _GEN_117;
  wire [26:0] _GEN_3330;
  wire [26:0] _T_7400;
  wire [26:0] _GEN_3331;
  wire [26:0] _T_7404;
  wire  _T_7424;
  wire  _GEN_118;
  wire [27:0] _GEN_3332;
  wire [27:0] _T_7440;
  wire [27:0] _GEN_3333;
  wire [27:0] _T_7444;
  wire  _T_7464;
  wire  _GEN_119;
  wire [28:0] _GEN_3334;
  wire [28:0] _T_7480;
  wire [28:0] _GEN_3335;
  wire [28:0] _T_7484;
  wire  _T_7504;
  wire  _GEN_120;
  wire [29:0] _GEN_3336;
  wire [29:0] _T_7520;
  wire [29:0] _GEN_3337;
  wire [29:0] _T_7524;
  wire  _T_7544;
  wire  _GEN_121;
  wire [30:0] _GEN_3338;
  wire [30:0] _T_7560;
  wire [30:0] _GEN_3339;
  wire [30:0] _T_7564;
  wire  _T_7584;
  wire  _GEN_122;
  wire [31:0] _GEN_3340;
  wire [31:0] _T_7600;
  wire [31:0] _GEN_3341;
  wire [31:0] _T_7604;
  wire  _T_7624;
  wire [31:0] _GEN_123;
  wire [31:0] _T_7643;
  wire  _T_7664;
  wire [31:0] _GEN_124;
  wire [31:0] _T_7683;
  wire  _T_7704;
  wire [31:0] _GEN_125;
  wire [31:0] _T_7723;
  wire  _T_7744;
  wire [31:0] _GEN_126;
  wire [31:0] _T_7763;
  wire  _T_7784;
  wire [31:0] _GEN_127;
  wire [31:0] _T_7803;
  wire  _T_7864;
  wire [31:0] _GEN_128;
  wire [31:0] _T_7883;
  wire  _T_7904;
  wire [31:0] _GEN_129;
  wire [31:0] _T_7923;
  wire  _T_7944;
  wire [31:0] _GEN_130;
  wire [31:0] _T_7963;
  wire  _T_7984;
  wire [31:0] _GEN_131;
  wire [31:0] _T_8003;
  wire  _T_8024;
  wire [31:0] _GEN_132;
  wire [31:0] _T_8043;
  wire  _T_8064;
  wire [31:0] _GEN_133;
  wire [31:0] _T_8083;
  wire  _T_8104;
  wire [31:0] _GEN_134;
  wire [31:0] _T_8123;
  wire  _T_8144;
  wire [31:0] _GEN_135;
  wire [31:0] _T_8163;
  wire  _T_8184;
  wire [31:0] _GEN_136;
  wire [31:0] _T_8203;
  wire  _T_8224;
  wire [31:0] _GEN_137;
  wire [31:0] _T_8243;
  wire  _T_8264;
  wire [31:0] _GEN_138;
  wire [31:0] _T_8283;
  wire  _T_8317;
  wire  _T_8318;
  wire  _T_8319;
  wire  _T_8320;
  wire  _T_8321;
  wire  _T_8322;
  wire  _T_8327;
  wire  _T_8328;
  wire  _T_8336;
  wire [1:0] _T_8341;
  wire [1:0] _T_8342;
  wire [3:0] _T_8343;
  wire [1:0] _T_8344;
  wire [1:0] _T_8345;
  wire [2:0] _T_8346;
  wire [4:0] _T_8347;
  wire [8:0] _T_8348;
  wire [511:0] _T_8864;
  wire  _T_8866;
  wire  _T_8867;
  wire  _T_8868;
  wire  _T_8869;
  wire  _T_8870;
  wire  _T_8871;
  wire  _T_8872;
  wire  _T_8873;
  wire  _T_8874;
  wire  _T_8875;
  wire  _T_8876;
  wire  _T_8877;
  wire  _T_8878;
  wire  _T_8879;
  wire  _T_8880;
  wire  _T_8881;
  wire  _T_8882;
  wire  _T_8883;
  wire  _T_8884;
  wire  _T_8885;
  wire  _T_8886;
  wire  _T_8887;
  wire  _T_8888;
  wire  _T_8889;
  wire  _T_8890;
  wire  _T_8891;
  wire  _T_8892;
  wire  _T_8893;
  wire  _T_8894;
  wire  _T_8895;
  wire  _T_8896;
  wire  _T_8897;
  wire  _T_8993;
  wire  _T_8994;
  wire  _T_9121;
  wire  _T_9122;
  wire  _T_18609;
  wire  _T_18610;
  wire  _T_20669;
  wire  _T_20670;
  wire  _T_23226;
  wire  _T_23227;
  wire  _T_23238;
  wire  _T_23239;
  wire  _T_23246;
  wire  _T_23247;
  wire  _T_23254;
  wire  _T_23255;
  wire  _T_23262;
  wire  _T_23263;
  wire  _T_23270;
  wire  _T_23271;
  wire  _T_23278;
  wire  _T_23279;
  wire  _T_23286;
  wire  _T_23287;
  wire  _T_23294;
  wire  _T_23295;
  wire  _T_23302;
  wire  _T_23303;
  wire  _T_23310;
  wire  _T_23311;
  wire  _T_23318;
  wire  _T_23319;
  wire  _T_23326;
  wire  _T_23327;
  wire  _T_23334;
  wire  _T_23335;
  wire  _T_23342;
  wire  _T_23343;
  wire  _T_23350;
  wire  _T_23351;
  wire  _T_23358;
  wire  _T_23359;
  wire  _T_23366;
  wire  _T_23367;
  wire  _T_23374;
  wire  _T_23375;
  wire  _T_23382;
  wire  _T_23383;
  wire  _T_23390;
  wire  _T_23391;
  wire  _T_23398;
  wire  _T_23399;
  wire  _T_23406;
  wire  _T_23407;
  wire  _T_23414;
  wire  _T_23415;
  wire  _T_23422;
  wire  _T_23423;
  wire  _T_23430;
  wire  _T_23431;
  wire  _T_23438;
  wire  _T_23439;
  wire  _T_23446;
  wire  _T_23447;
  wire  _T_23454;
  wire  _T_23455;
  wire  _T_23462;
  wire  _T_23463;
  wire  _T_23470;
  wire  _T_23471;
  wire  _T_23478;
  wire  _T_23479;
  wire  _T_23486;
  wire  _T_23487;
  wire  _T_24254;
  wire  _T_24255;
  wire  _T_24262;
  wire  _T_24263;
  wire  _T_25278;
  wire  _T_25279;
  wire  _T_25286;
  wire  _T_25287;
  wire  _T_27850;
  wire  _T_27853_0;
  wire  _T_27853_1;
  wire  _T_27853_2;
  wire  _T_27853_3;
  wire  _T_27853_4;
  wire  _T_27853_5;
  wire  _T_27853_6;
  wire  _T_27853_7;
  wire  _T_27853_8;
  wire  _T_27853_9;
  wire  _T_27853_10;
  wire  _T_27853_11;
  wire  _T_27853_12;
  wire  _T_27853_13;
  wire  _T_27853_14;
  wire  _T_27853_15;
  wire  _T_27853_16;
  wire  _T_27853_17;
  wire  _T_27853_18;
  wire  _T_27853_19;
  wire  _T_27853_20;
  wire  _T_27853_21;
  wire  _T_27853_22;
  wire  _T_27853_23;
  wire  _T_27853_24;
  wire  _T_27853_25;
  wire  _T_27853_26;
  wire  _T_27853_27;
  wire  _T_27853_28;
  wire  _T_27853_29;
  wire  _T_27853_30;
  wire  _T_27853_31;
  wire  _T_27853_32;
  wire  _T_27853_64;
  wire  _T_27853_65;
  wire  _T_27853_128;
  wire  _T_27853_129;
  wire  _T_27853_256;
  wire  _T_27853_257;
  wire [31:0] _T_28371_1;
  wire [31:0] _T_28371_2;
  wire [31:0] _T_28371_3;
  wire [31:0] _T_28371_4;
  wire [31:0] _T_28371_5;
  wire [31:0] _T_28371_6;
  wire [31:0] _T_28371_7;
  wire [31:0] _T_28371_8;
  wire [31:0] _T_28371_9;
  wire [31:0] _T_28371_10;
  wire [31:0] _T_28371_11;
  wire [31:0] _T_28371_12;
  wire [31:0] _T_28371_13;
  wire [31:0] _T_28371_14;
  wire [31:0] _T_28371_15;
  wire [31:0] _T_28371_16;
  wire [31:0] _T_28371_17;
  wire [31:0] _T_28371_18;
  wire [31:0] _T_28371_19;
  wire [31:0] _T_28371_20;
  wire [31:0] _T_28371_21;
  wire [31:0] _T_28371_22;
  wire [31:0] _T_28371_23;
  wire [31:0] _T_28371_24;
  wire [31:0] _T_28371_25;
  wire [31:0] _T_28371_26;
  wire [31:0] _T_28371_27;
  wire [31:0] _T_28371_28;
  wire [31:0] _T_28371_29;
  wire [31:0] _T_28371_30;
  wire [31:0] _T_28371_31;
  wire [31:0] _T_28371_32;
  wire [31:0] _T_28371_64;
  wire [31:0] _T_28371_65;
  wire [31:0] _T_28371_128;
  wire [31:0] _T_28371_129;
  wire [31:0] _T_28371_256;
  wire [31:0] _T_28371_257;
  wire  _GEN_5;
  wire  _GEN_2183;
  wire  _GEN_2184;
  wire  _GEN_2185;
  wire  _GEN_2186;
  wire  _GEN_2187;
  wire  _GEN_2188;
  wire  _GEN_2189;
  wire  _GEN_2190;
  wire  _GEN_2191;
  wire  _GEN_2192;
  wire  _GEN_2193;
  wire  _GEN_2194;
  wire  _GEN_2195;
  wire  _GEN_2196;
  wire  _GEN_2197;
  wire  _GEN_2198;
  wire  _GEN_2199;
  wire  _GEN_2200;
  wire  _GEN_2201;
  wire  _GEN_2202;
  wire  _GEN_2203;
  wire  _GEN_2204;
  wire  _GEN_2205;
  wire  _GEN_2206;
  wire  _GEN_2207;
  wire  _GEN_2208;
  wire  _GEN_2209;
  wire  _GEN_2210;
  wire  _GEN_2211;
  wire  _GEN_2212;
  wire  _GEN_2213;
  wire  _GEN_2214;
  wire  _GEN_2215;
  wire  _GEN_2216;
  wire  _GEN_2217;
  wire  _GEN_2218;
  wire  _GEN_2219;
  wire  _GEN_2220;
  wire  _GEN_2221;
  wire  _GEN_2222;
  wire  _GEN_2223;
  wire  _GEN_2224;
  wire  _GEN_2225;
  wire  _GEN_2226;
  wire  _GEN_2227;
  wire  _GEN_2228;
  wire  _GEN_2229;
  wire  _GEN_2230;
  wire  _GEN_2231;
  wire  _GEN_2232;
  wire  _GEN_2233;
  wire  _GEN_2234;
  wire  _GEN_2235;
  wire  _GEN_2236;
  wire  _GEN_2237;
  wire  _GEN_2238;
  wire  _GEN_2239;
  wire  _GEN_2240;
  wire  _GEN_2241;
  wire  _GEN_2242;
  wire  _GEN_2243;
  wire  _GEN_2244;
  wire  _GEN_2245;
  wire  _GEN_2246;
  wire  _GEN_2247;
  wire  _GEN_2248;
  wire  _GEN_2249;
  wire  _GEN_2250;
  wire  _GEN_2251;
  wire  _GEN_2252;
  wire  _GEN_2253;
  wire  _GEN_2254;
  wire  _GEN_2255;
  wire  _GEN_2256;
  wire  _GEN_2257;
  wire  _GEN_2258;
  wire  _GEN_2259;
  wire  _GEN_2260;
  wire  _GEN_2261;
  wire  _GEN_2262;
  wire  _GEN_2263;
  wire  _GEN_2264;
  wire  _GEN_2265;
  wire  _GEN_2266;
  wire  _GEN_2267;
  wire  _GEN_2268;
  wire  _GEN_2269;
  wire  _GEN_2270;
  wire  _GEN_2271;
  wire  _GEN_2272;
  wire  _GEN_2273;
  wire  _GEN_2274;
  wire  _GEN_2275;
  wire  _GEN_2276;
  wire  _GEN_2277;
  wire  _GEN_2278;
  wire  _GEN_2279;
  wire  _GEN_2280;
  wire  _GEN_2281;
  wire  _GEN_2282;
  wire  _GEN_2283;
  wire  _GEN_2284;
  wire  _GEN_2285;
  wire  _GEN_2286;
  wire  _GEN_2287;
  wire  _GEN_2288;
  wire  _GEN_2289;
  wire  _GEN_2290;
  wire  _GEN_2291;
  wire  _GEN_2292;
  wire  _GEN_2293;
  wire  _GEN_2294;
  wire  _GEN_2295;
  wire  _GEN_2296;
  wire  _GEN_2297;
  wire  _GEN_2298;
  wire  _GEN_2299;
  wire  _GEN_2300;
  wire  _GEN_2301;
  wire  _GEN_2302;
  wire  _GEN_2303;
  wire  _GEN_2304;
  wire  _GEN_2305;
  wire  _GEN_2306;
  wire  _GEN_2307;
  wire  _GEN_2308;
  wire  _GEN_2309;
  wire  _GEN_2310;
  wire  _GEN_2311;
  wire  _GEN_2312;
  wire  _GEN_2313;
  wire  _GEN_2314;
  wire  _GEN_2315;
  wire  _GEN_2316;
  wire  _GEN_2317;
  wire  _GEN_2318;
  wire  _GEN_2319;
  wire  _GEN_2320;
  wire  _GEN_2321;
  wire  _GEN_2322;
  wire  _GEN_2323;
  wire  _GEN_2324;
  wire  _GEN_2325;
  wire  _GEN_2326;
  wire  _GEN_2327;
  wire  _GEN_2328;
  wire  _GEN_2329;
  wire  _GEN_2330;
  wire  _GEN_2331;
  wire  _GEN_2332;
  wire  _GEN_2333;
  wire  _GEN_2334;
  wire  _GEN_2335;
  wire  _GEN_2336;
  wire  _GEN_2337;
  wire  _GEN_2338;
  wire  _GEN_2339;
  wire  _GEN_2340;
  wire  _GEN_2341;
  wire  _GEN_2342;
  wire  _GEN_2343;
  wire  _GEN_2344;
  wire  _GEN_2345;
  wire  _GEN_2346;
  wire  _GEN_2347;
  wire  _GEN_2348;
  wire  _GEN_2349;
  wire  _GEN_2350;
  wire  _GEN_2351;
  wire  _GEN_2352;
  wire  _GEN_2353;
  wire  _GEN_2354;
  wire  _GEN_2355;
  wire  _GEN_2356;
  wire  _GEN_2357;
  wire  _GEN_2358;
  wire  _GEN_2359;
  wire  _GEN_2360;
  wire  _GEN_2361;
  wire  _GEN_2362;
  wire  _GEN_2363;
  wire  _GEN_2364;
  wire  _GEN_2365;
  wire  _GEN_2366;
  wire  _GEN_2367;
  wire  _GEN_2368;
  wire  _GEN_2369;
  wire  _GEN_2370;
  wire  _GEN_2371;
  wire  _GEN_2372;
  wire  _GEN_2373;
  wire  _GEN_2374;
  wire  _GEN_2375;
  wire  _GEN_2376;
  wire  _GEN_2377;
  wire  _GEN_2378;
  wire  _GEN_2379;
  wire  _GEN_2380;
  wire  _GEN_2381;
  wire  _GEN_2382;
  wire  _GEN_2383;
  wire  _GEN_2384;
  wire  _GEN_2385;
  wire  _GEN_2386;
  wire  _GEN_2387;
  wire  _GEN_2388;
  wire  _GEN_2389;
  wire  _GEN_2390;
  wire  _GEN_2391;
  wire  _GEN_2392;
  wire  _GEN_2393;
  wire  _GEN_2394;
  wire  _GEN_2395;
  wire  _GEN_2396;
  wire  _GEN_2397;
  wire  _GEN_2398;
  wire  _GEN_2399;
  wire  _GEN_2400;
  wire  _GEN_2401;
  wire  _GEN_2402;
  wire  _GEN_2403;
  wire  _GEN_2404;
  wire  _GEN_2405;
  wire  _GEN_2406;
  wire  _GEN_2407;
  wire  _GEN_2408;
  wire  _GEN_2409;
  wire  _GEN_2410;
  wire  _GEN_2411;
  wire  _GEN_2412;
  wire  _GEN_2413;
  wire  _GEN_2414;
  wire  _GEN_2415;
  wire  _GEN_2416;
  wire  _GEN_2417;
  wire  _GEN_2418;
  wire  _GEN_2419;
  wire  _GEN_2420;
  wire  _GEN_2421;
  wire  _GEN_2422;
  wire  _GEN_2423;
  wire  _GEN_2424;
  wire  _GEN_2425;
  wire  _GEN_2426;
  wire  _GEN_2427;
  wire  _GEN_2428;
  wire  _GEN_2429;
  wire  _GEN_2430;
  wire  _GEN_2431;
  wire  _GEN_2432;
  wire  _GEN_2433;
  wire  _GEN_2434;
  wire  _GEN_2435;
  wire  _GEN_2436;
  wire  _GEN_2437;
  wire  _GEN_2438;
  wire  _GEN_2439;
  wire  _GEN_2440;
  wire  _GEN_2441;
  wire  _GEN_2442;
  wire  _GEN_2443;
  wire  _GEN_2444;
  wire  _GEN_2445;
  wire  _GEN_2446;
  wire  _GEN_2447;
  wire  _GEN_2448;
  wire  _GEN_2449;
  wire  _GEN_2450;
  wire  _GEN_2451;
  wire  _GEN_2452;
  wire  _GEN_2453;
  wire  _GEN_2454;
  wire  _GEN_2455;
  wire  _GEN_2456;
  wire  _GEN_2457;
  wire  _GEN_2458;
  wire  _GEN_2459;
  wire  _GEN_2460;
  wire  _GEN_2461;
  wire  _GEN_2462;
  wire  _GEN_2463;
  wire  _GEN_2464;
  wire  _GEN_2465;
  wire  _GEN_2466;
  wire  _GEN_2467;
  wire  _GEN_2468;
  wire  _GEN_2469;
  wire  _GEN_2470;
  wire  _GEN_2471;
  wire  _GEN_2472;
  wire  _GEN_2473;
  wire  _GEN_2474;
  wire  _GEN_2475;
  wire  _GEN_2476;
  wire  _GEN_2477;
  wire  _GEN_2478;
  wire  _GEN_2479;
  wire  _GEN_2480;
  wire  _GEN_2481;
  wire  _GEN_2482;
  wire  _GEN_2483;
  wire  _GEN_2484;
  wire  _GEN_2485;
  wire  _GEN_2486;
  wire  _GEN_2487;
  wire  _GEN_2488;
  wire  _GEN_2489;
  wire  _GEN_2490;
  wire  _GEN_2491;
  wire  _GEN_2492;
  wire  _GEN_2493;
  wire  _GEN_2494;
  wire  _GEN_2495;
  wire  _GEN_2496;
  wire  _GEN_2497;
  wire  _GEN_2498;
  wire  _GEN_2499;
  wire  _GEN_2500;
  wire  _GEN_2501;
  wire  _GEN_2502;
  wire  _GEN_2503;
  wire  _GEN_2504;
  wire  _GEN_2505;
  wire  _GEN_2506;
  wire  _GEN_2507;
  wire  _GEN_2508;
  wire  _GEN_2509;
  wire  _GEN_2510;
  wire  _GEN_2511;
  wire  _GEN_2512;
  wire  _GEN_2513;
  wire  _GEN_2514;
  wire  _GEN_2515;
  wire  _GEN_2516;
  wire  _GEN_2517;
  wire  _GEN_2518;
  wire  _GEN_2519;
  wire  _GEN_2520;
  wire  _GEN_2521;
  wire  _GEN_2522;
  wire  _GEN_2523;
  wire  _GEN_2524;
  wire  _GEN_2525;
  wire  _GEN_2526;
  wire  _GEN_2527;
  wire  _GEN_2528;
  wire  _GEN_2529;
  wire  _GEN_2530;
  wire  _GEN_2531;
  wire  _GEN_2532;
  wire  _GEN_2533;
  wire  _GEN_2534;
  wire  _GEN_2535;
  wire  _GEN_2536;
  wire  _GEN_2537;
  wire  _GEN_2538;
  wire  _GEN_2539;
  wire  _GEN_2540;
  wire  _GEN_2541;
  wire  _GEN_2542;
  wire  _GEN_2543;
  wire  _GEN_2544;
  wire  _GEN_2545;
  wire  _GEN_2546;
  wire  _GEN_2547;
  wire  _GEN_2548;
  wire  _GEN_2549;
  wire  _GEN_2550;
  wire  _GEN_2551;
  wire  _GEN_2552;
  wire  _GEN_2553;
  wire  _GEN_2554;
  wire  _GEN_2555;
  wire  _GEN_2556;
  wire  _GEN_2557;
  wire  _GEN_2558;
  wire  _GEN_2559;
  wire  _GEN_2560;
  wire  _GEN_2561;
  wire  _GEN_2562;
  wire  _GEN_2563;
  wire  _GEN_2564;
  wire  _GEN_2565;
  wire  _GEN_2566;
  wire  _GEN_2567;
  wire  _GEN_2568;
  wire  _GEN_2569;
  wire  _GEN_2570;
  wire  _GEN_2571;
  wire  _GEN_2572;
  wire  _GEN_2573;
  wire  _GEN_2574;
  wire  _GEN_2575;
  wire  _GEN_2576;
  wire  _GEN_2577;
  wire  _GEN_2578;
  wire  _GEN_2579;
  wire  _GEN_2580;
  wire  _GEN_2581;
  wire  _GEN_2582;
  wire  _GEN_2583;
  wire  _GEN_2584;
  wire  _GEN_2585;
  wire  _GEN_2586;
  wire  _GEN_2587;
  wire  _GEN_2588;
  wire  _GEN_2589;
  wire  _GEN_2590;
  wire  _GEN_2591;
  wire  _GEN_2592;
  wire  _GEN_2593;
  wire  _GEN_2594;
  wire  _GEN_2595;
  wire  _GEN_2596;
  wire  _GEN_2597;
  wire  _GEN_2598;
  wire  _GEN_2599;
  wire  _GEN_2600;
  wire  _GEN_2601;
  wire  _GEN_2602;
  wire  _GEN_2603;
  wire  _GEN_2604;
  wire  _GEN_2605;
  wire  _GEN_2606;
  wire  _GEN_2607;
  wire  _GEN_2608;
  wire  _GEN_2609;
  wire  _GEN_2610;
  wire  _GEN_2611;
  wire  _GEN_2612;
  wire  _GEN_2613;
  wire  _GEN_2614;
  wire  _GEN_2615;
  wire  _GEN_2616;
  wire  _GEN_2617;
  wire  _GEN_2618;
  wire  _GEN_2619;
  wire  _GEN_2620;
  wire  _GEN_2621;
  wire  _GEN_2622;
  wire  _GEN_2623;
  wire  _GEN_2624;
  wire  _GEN_2625;
  wire  _GEN_2626;
  wire  _GEN_2627;
  wire  _GEN_2628;
  wire  _GEN_2629;
  wire  _GEN_2630;
  wire  _GEN_2631;
  wire  _GEN_2632;
  wire  _GEN_2633;
  wire  _GEN_2634;
  wire  _GEN_2635;
  wire  _GEN_2636;
  wire  _GEN_2637;
  wire  _GEN_2638;
  wire  _GEN_2639;
  wire  _GEN_2640;
  wire  _GEN_2641;
  wire  _GEN_2642;
  wire  _GEN_2643;
  wire  _GEN_2644;
  wire  _GEN_2645;
  wire  _GEN_2646;
  wire  _GEN_2647;
  wire  _GEN_2648;
  wire  _GEN_2649;
  wire  _GEN_2650;
  wire  _GEN_2651;
  wire  _GEN_2652;
  wire  _GEN_2653;
  wire  _GEN_2654;
  wire  _GEN_2655;
  wire  _GEN_2656;
  wire  _GEN_2657;
  wire  _GEN_2658;
  wire  _GEN_2659;
  wire  _GEN_2660;
  wire  _GEN_2661;
  wire  _GEN_2662;
  wire  _GEN_2663;
  wire  _GEN_2664;
  wire  _GEN_2665;
  wire  _GEN_2666;
  wire  _GEN_2667;
  wire  _GEN_2668;
  wire  _GEN_2669;
  wire  _GEN_2670;
  wire  _GEN_2671;
  wire  _GEN_2672;
  wire  _GEN_2673;
  wire  _GEN_2674;
  wire  _GEN_2675;
  wire  _GEN_2676;
  wire  _GEN_2677;
  wire  _GEN_2678;
  wire  _GEN_2679;
  wire  _GEN_2680;
  wire  _GEN_2681;
  wire  _GEN_2682;
  wire  _GEN_2683;
  wire  _GEN_2684;
  wire  _GEN_2685;
  wire  _GEN_2686;
  wire  _GEN_2687;
  wire  _GEN_2688;
  wire  _GEN_2689;
  wire  _GEN_2690;
  wire  _GEN_2691;
  wire  _GEN_2692;
  wire  _GEN_2693;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_2694;
  wire [31:0] _GEN_2695;
  wire [31:0] _GEN_2696;
  wire [31:0] _GEN_2697;
  wire [31:0] _GEN_2698;
  wire [31:0] _GEN_2699;
  wire [31:0] _GEN_2700;
  wire [31:0] _GEN_2701;
  wire [31:0] _GEN_2702;
  wire [31:0] _GEN_2703;
  wire [31:0] _GEN_2704;
  wire [31:0] _GEN_2705;
  wire [31:0] _GEN_2706;
  wire [31:0] _GEN_2707;
  wire [31:0] _GEN_2708;
  wire [31:0] _GEN_2709;
  wire [31:0] _GEN_2710;
  wire [31:0] _GEN_2711;
  wire [31:0] _GEN_2712;
  wire [31:0] _GEN_2713;
  wire [31:0] _GEN_2714;
  wire [31:0] _GEN_2715;
  wire [31:0] _GEN_2716;
  wire [31:0] _GEN_2717;
  wire [31:0] _GEN_2718;
  wire [31:0] _GEN_2719;
  wire [31:0] _GEN_2720;
  wire [31:0] _GEN_2721;
  wire [31:0] _GEN_2722;
  wire [31:0] _GEN_2723;
  wire [31:0] _GEN_2724;
  wire [31:0] _GEN_2725;
  wire [31:0] _GEN_2726;
  wire [31:0] _GEN_2727;
  wire [31:0] _GEN_2728;
  wire [31:0] _GEN_2729;
  wire [31:0] _GEN_2730;
  wire [31:0] _GEN_2731;
  wire [31:0] _GEN_2732;
  wire [31:0] _GEN_2733;
  wire [31:0] _GEN_2734;
  wire [31:0] _GEN_2735;
  wire [31:0] _GEN_2736;
  wire [31:0] _GEN_2737;
  wire [31:0] _GEN_2738;
  wire [31:0] _GEN_2739;
  wire [31:0] _GEN_2740;
  wire [31:0] _GEN_2741;
  wire [31:0] _GEN_2742;
  wire [31:0] _GEN_2743;
  wire [31:0] _GEN_2744;
  wire [31:0] _GEN_2745;
  wire [31:0] _GEN_2746;
  wire [31:0] _GEN_2747;
  wire [31:0] _GEN_2748;
  wire [31:0] _GEN_2749;
  wire [31:0] _GEN_2750;
  wire [31:0] _GEN_2751;
  wire [31:0] _GEN_2752;
  wire [31:0] _GEN_2753;
  wire [31:0] _GEN_2754;
  wire [31:0] _GEN_2755;
  wire [31:0] _GEN_2756;
  wire [31:0] _GEN_2757;
  wire [31:0] _GEN_2758;
  wire [31:0] _GEN_2759;
  wire [31:0] _GEN_2760;
  wire [31:0] _GEN_2761;
  wire [31:0] _GEN_2762;
  wire [31:0] _GEN_2763;
  wire [31:0] _GEN_2764;
  wire [31:0] _GEN_2765;
  wire [31:0] _GEN_2766;
  wire [31:0] _GEN_2767;
  wire [31:0] _GEN_2768;
  wire [31:0] _GEN_2769;
  wire [31:0] _GEN_2770;
  wire [31:0] _GEN_2771;
  wire [31:0] _GEN_2772;
  wire [31:0] _GEN_2773;
  wire [31:0] _GEN_2774;
  wire [31:0] _GEN_2775;
  wire [31:0] _GEN_2776;
  wire [31:0] _GEN_2777;
  wire [31:0] _GEN_2778;
  wire [31:0] _GEN_2779;
  wire [31:0] _GEN_2780;
  wire [31:0] _GEN_2781;
  wire [31:0] _GEN_2782;
  wire [31:0] _GEN_2783;
  wire [31:0] _GEN_2784;
  wire [31:0] _GEN_2785;
  wire [31:0] _GEN_2786;
  wire [31:0] _GEN_2787;
  wire [31:0] _GEN_2788;
  wire [31:0] _GEN_2789;
  wire [31:0] _GEN_2790;
  wire [31:0] _GEN_2791;
  wire [31:0] _GEN_2792;
  wire [31:0] _GEN_2793;
  wire [31:0] _GEN_2794;
  wire [31:0] _GEN_2795;
  wire [31:0] _GEN_2796;
  wire [31:0] _GEN_2797;
  wire [31:0] _GEN_2798;
  wire [31:0] _GEN_2799;
  wire [31:0] _GEN_2800;
  wire [31:0] _GEN_2801;
  wire [31:0] _GEN_2802;
  wire [31:0] _GEN_2803;
  wire [31:0] _GEN_2804;
  wire [31:0] _GEN_2805;
  wire [31:0] _GEN_2806;
  wire [31:0] _GEN_2807;
  wire [31:0] _GEN_2808;
  wire [31:0] _GEN_2809;
  wire [31:0] _GEN_2810;
  wire [31:0] _GEN_2811;
  wire [31:0] _GEN_2812;
  wire [31:0] _GEN_2813;
  wire [31:0] _GEN_2814;
  wire [31:0] _GEN_2815;
  wire [31:0] _GEN_2816;
  wire [31:0] _GEN_2817;
  wire [31:0] _GEN_2818;
  wire [31:0] _GEN_2819;
  wire [31:0] _GEN_2820;
  wire [31:0] _GEN_2821;
  wire [31:0] _GEN_2822;
  wire [31:0] _GEN_2823;
  wire [31:0] _GEN_2824;
  wire [31:0] _GEN_2825;
  wire [31:0] _GEN_2826;
  wire [31:0] _GEN_2827;
  wire [31:0] _GEN_2828;
  wire [31:0] _GEN_2829;
  wire [31:0] _GEN_2830;
  wire [31:0] _GEN_2831;
  wire [31:0] _GEN_2832;
  wire [31:0] _GEN_2833;
  wire [31:0] _GEN_2834;
  wire [31:0] _GEN_2835;
  wire [31:0] _GEN_2836;
  wire [31:0] _GEN_2837;
  wire [31:0] _GEN_2838;
  wire [31:0] _GEN_2839;
  wire [31:0] _GEN_2840;
  wire [31:0] _GEN_2841;
  wire [31:0] _GEN_2842;
  wire [31:0] _GEN_2843;
  wire [31:0] _GEN_2844;
  wire [31:0] _GEN_2845;
  wire [31:0] _GEN_2846;
  wire [31:0] _GEN_2847;
  wire [31:0] _GEN_2848;
  wire [31:0] _GEN_2849;
  wire [31:0] _GEN_2850;
  wire [31:0] _GEN_2851;
  wire [31:0] _GEN_2852;
  wire [31:0] _GEN_2853;
  wire [31:0] _GEN_2854;
  wire [31:0] _GEN_2855;
  wire [31:0] _GEN_2856;
  wire [31:0] _GEN_2857;
  wire [31:0] _GEN_2858;
  wire [31:0] _GEN_2859;
  wire [31:0] _GEN_2860;
  wire [31:0] _GEN_2861;
  wire [31:0] _GEN_2862;
  wire [31:0] _GEN_2863;
  wire [31:0] _GEN_2864;
  wire [31:0] _GEN_2865;
  wire [31:0] _GEN_2866;
  wire [31:0] _GEN_2867;
  wire [31:0] _GEN_2868;
  wire [31:0] _GEN_2869;
  wire [31:0] _GEN_2870;
  wire [31:0] _GEN_2871;
  wire [31:0] _GEN_2872;
  wire [31:0] _GEN_2873;
  wire [31:0] _GEN_2874;
  wire [31:0] _GEN_2875;
  wire [31:0] _GEN_2876;
  wire [31:0] _GEN_2877;
  wire [31:0] _GEN_2878;
  wire [31:0] _GEN_2879;
  wire [31:0] _GEN_2880;
  wire [31:0] _GEN_2881;
  wire [31:0] _GEN_2882;
  wire [31:0] _GEN_2883;
  wire [31:0] _GEN_2884;
  wire [31:0] _GEN_2885;
  wire [31:0] _GEN_2886;
  wire [31:0] _GEN_2887;
  wire [31:0] _GEN_2888;
  wire [31:0] _GEN_2889;
  wire [31:0] _GEN_2890;
  wire [31:0] _GEN_2891;
  wire [31:0] _GEN_2892;
  wire [31:0] _GEN_2893;
  wire [31:0] _GEN_2894;
  wire [31:0] _GEN_2895;
  wire [31:0] _GEN_2896;
  wire [31:0] _GEN_2897;
  wire [31:0] _GEN_2898;
  wire [31:0] _GEN_2899;
  wire [31:0] _GEN_2900;
  wire [31:0] _GEN_2901;
  wire [31:0] _GEN_2902;
  wire [31:0] _GEN_2903;
  wire [31:0] _GEN_2904;
  wire [31:0] _GEN_2905;
  wire [31:0] _GEN_2906;
  wire [31:0] _GEN_2907;
  wire [31:0] _GEN_2908;
  wire [31:0] _GEN_2909;
  wire [31:0] _GEN_2910;
  wire [31:0] _GEN_2911;
  wire [31:0] _GEN_2912;
  wire [31:0] _GEN_2913;
  wire [31:0] _GEN_2914;
  wire [31:0] _GEN_2915;
  wire [31:0] _GEN_2916;
  wire [31:0] _GEN_2917;
  wire [31:0] _GEN_2918;
  wire [31:0] _GEN_2919;
  wire [31:0] _GEN_2920;
  wire [31:0] _GEN_2921;
  wire [31:0] _GEN_2922;
  wire [31:0] _GEN_2923;
  wire [31:0] _GEN_2924;
  wire [31:0] _GEN_2925;
  wire [31:0] _GEN_2926;
  wire [31:0] _GEN_2927;
  wire [31:0] _GEN_2928;
  wire [31:0] _GEN_2929;
  wire [31:0] _GEN_2930;
  wire [31:0] _GEN_2931;
  wire [31:0] _GEN_2932;
  wire [31:0] _GEN_2933;
  wire [31:0] _GEN_2934;
  wire [31:0] _GEN_2935;
  wire [31:0] _GEN_2936;
  wire [31:0] _GEN_2937;
  wire [31:0] _GEN_2938;
  wire [31:0] _GEN_2939;
  wire [31:0] _GEN_2940;
  wire [31:0] _GEN_2941;
  wire [31:0] _GEN_2942;
  wire [31:0] _GEN_2943;
  wire [31:0] _GEN_2944;
  wire [31:0] _GEN_2945;
  wire [31:0] _GEN_2946;
  wire [31:0] _GEN_2947;
  wire [31:0] _GEN_2948;
  wire [31:0] _GEN_2949;
  wire [31:0] _GEN_2950;
  wire [31:0] _GEN_2951;
  wire [31:0] _GEN_2952;
  wire [31:0] _GEN_2953;
  wire [31:0] _GEN_2954;
  wire [31:0] _GEN_2955;
  wire [31:0] _GEN_2956;
  wire [31:0] _GEN_2957;
  wire [31:0] _GEN_2958;
  wire [31:0] _GEN_2959;
  wire [31:0] _GEN_2960;
  wire [31:0] _GEN_2961;
  wire [31:0] _GEN_2962;
  wire [31:0] _GEN_2963;
  wire [31:0] _GEN_2964;
  wire [31:0] _GEN_2965;
  wire [31:0] _GEN_2966;
  wire [31:0] _GEN_2967;
  wire [31:0] _GEN_2968;
  wire [31:0] _GEN_2969;
  wire [31:0] _GEN_2970;
  wire [31:0] _GEN_2971;
  wire [31:0] _GEN_2972;
  wire [31:0] _GEN_2973;
  wire [31:0] _GEN_2974;
  wire [31:0] _GEN_2975;
  wire [31:0] _GEN_2976;
  wire [31:0] _GEN_2977;
  wire [31:0] _GEN_2978;
  wire [31:0] _GEN_2979;
  wire [31:0] _GEN_2980;
  wire [31:0] _GEN_2981;
  wire [31:0] _GEN_2982;
  wire [31:0] _GEN_2983;
  wire [31:0] _GEN_2984;
  wire [31:0] _GEN_2985;
  wire [31:0] _GEN_2986;
  wire [31:0] _GEN_2987;
  wire [31:0] _GEN_2988;
  wire [31:0] _GEN_2989;
  wire [31:0] _GEN_2990;
  wire [31:0] _GEN_2991;
  wire [31:0] _GEN_2992;
  wire [31:0] _GEN_2993;
  wire [31:0] _GEN_2994;
  wire [31:0] _GEN_2995;
  wire [31:0] _GEN_2996;
  wire [31:0] _GEN_2997;
  wire [31:0] _GEN_2998;
  wire [31:0] _GEN_2999;
  wire [31:0] _GEN_3000;
  wire [31:0] _GEN_3001;
  wire [31:0] _GEN_3002;
  wire [31:0] _GEN_3003;
  wire [31:0] _GEN_3004;
  wire [31:0] _GEN_3005;
  wire [31:0] _GEN_3006;
  wire [31:0] _GEN_3007;
  wire [31:0] _GEN_3008;
  wire [31:0] _GEN_3009;
  wire [31:0] _GEN_3010;
  wire [31:0] _GEN_3011;
  wire [31:0] _GEN_3012;
  wire [31:0] _GEN_3013;
  wire [31:0] _GEN_3014;
  wire [31:0] _GEN_3015;
  wire [31:0] _GEN_3016;
  wire [31:0] _GEN_3017;
  wire [31:0] _GEN_3018;
  wire [31:0] _GEN_3019;
  wire [31:0] _GEN_3020;
  wire [31:0] _GEN_3021;
  wire [31:0] _GEN_3022;
  wire [31:0] _GEN_3023;
  wire [31:0] _GEN_3024;
  wire [31:0] _GEN_3025;
  wire [31:0] _GEN_3026;
  wire [31:0] _GEN_3027;
  wire [31:0] _GEN_3028;
  wire [31:0] _GEN_3029;
  wire [31:0] _GEN_3030;
  wire [31:0] _GEN_3031;
  wire [31:0] _GEN_3032;
  wire [31:0] _GEN_3033;
  wire [31:0] _GEN_3034;
  wire [31:0] _GEN_3035;
  wire [31:0] _GEN_3036;
  wire [31:0] _GEN_3037;
  wire [31:0] _GEN_3038;
  wire [31:0] _GEN_3039;
  wire [31:0] _GEN_3040;
  wire [31:0] _GEN_3041;
  wire [31:0] _GEN_3042;
  wire [31:0] _GEN_3043;
  wire [31:0] _GEN_3044;
  wire [31:0] _GEN_3045;
  wire [31:0] _GEN_3046;
  wire [31:0] _GEN_3047;
  wire [31:0] _GEN_3048;
  wire [31:0] _GEN_3049;
  wire [31:0] _GEN_3050;
  wire [31:0] _GEN_3051;
  wire [31:0] _GEN_3052;
  wire [31:0] _GEN_3053;
  wire [31:0] _GEN_3054;
  wire [31:0] _GEN_3055;
  wire [31:0] _GEN_3056;
  wire [31:0] _GEN_3057;
  wire [31:0] _GEN_3058;
  wire [31:0] _GEN_3059;
  wire [31:0] _GEN_3060;
  wire [31:0] _GEN_3061;
  wire [31:0] _GEN_3062;
  wire [31:0] _GEN_3063;
  wire [31:0] _GEN_3064;
  wire [31:0] _GEN_3065;
  wire [31:0] _GEN_3066;
  wire [31:0] _GEN_3067;
  wire [31:0] _GEN_3068;
  wire [31:0] _GEN_3069;
  wire [31:0] _GEN_3070;
  wire [31:0] _GEN_3071;
  wire [31:0] _GEN_3072;
  wire [31:0] _GEN_3073;
  wire [31:0] _GEN_3074;
  wire [31:0] _GEN_3075;
  wire [31:0] _GEN_3076;
  wire [31:0] _GEN_3077;
  wire [31:0] _GEN_3078;
  wire [31:0] _GEN_3079;
  wire [31:0] _GEN_3080;
  wire [31:0] _GEN_3081;
  wire [31:0] _GEN_3082;
  wire [31:0] _GEN_3083;
  wire [31:0] _GEN_3084;
  wire [31:0] _GEN_3085;
  wire [31:0] _GEN_3086;
  wire [31:0] _GEN_3087;
  wire [31:0] _GEN_3088;
  wire [31:0] _GEN_3089;
  wire [31:0] _GEN_3090;
  wire [31:0] _GEN_3091;
  wire [31:0] _GEN_3092;
  wire [31:0] _GEN_3093;
  wire [31:0] _GEN_3094;
  wire [31:0] _GEN_3095;
  wire [31:0] _GEN_3096;
  wire [31:0] _GEN_3097;
  wire [31:0] _GEN_3098;
  wire [31:0] _GEN_3099;
  wire [31:0] _GEN_3100;
  wire [31:0] _GEN_3101;
  wire [31:0] _GEN_3102;
  wire [31:0] _GEN_3103;
  wire [31:0] _GEN_3104;
  wire [31:0] _GEN_3105;
  wire [31:0] _GEN_3106;
  wire [31:0] _GEN_3107;
  wire [31:0] _GEN_3108;
  wire [31:0] _GEN_3109;
  wire [31:0] _GEN_3110;
  wire [31:0] _GEN_3111;
  wire [31:0] _GEN_3112;
  wire [31:0] _GEN_3113;
  wire [31:0] _GEN_3114;
  wire [31:0] _GEN_3115;
  wire [31:0] _GEN_3116;
  wire [31:0] _GEN_3117;
  wire [31:0] _GEN_3118;
  wire [31:0] _GEN_3119;
  wire [31:0] _GEN_3120;
  wire [31:0] _GEN_3121;
  wire [31:0] _GEN_3122;
  wire [31:0] _GEN_3123;
  wire [31:0] _GEN_3124;
  wire [31:0] _GEN_3125;
  wire [31:0] _GEN_3126;
  wire [31:0] _GEN_3127;
  wire [31:0] _GEN_3128;
  wire [31:0] _GEN_3129;
  wire [31:0] _GEN_3130;
  wire [31:0] _GEN_3131;
  wire [31:0] _GEN_3132;
  wire [31:0] _GEN_3133;
  wire [31:0] _GEN_3134;
  wire [31:0] _GEN_3135;
  wire [31:0] _GEN_3136;
  wire [31:0] _GEN_3137;
  wire [31:0] _GEN_3138;
  wire [31:0] _GEN_3139;
  wire [31:0] _GEN_3140;
  wire [31:0] _GEN_3141;
  wire [31:0] _GEN_3142;
  wire [31:0] _GEN_3143;
  wire [31:0] _GEN_3144;
  wire [31:0] _GEN_3145;
  wire [31:0] _GEN_3146;
  wire [31:0] _GEN_3147;
  wire [31:0] _GEN_3148;
  wire [31:0] _GEN_3149;
  wire [31:0] _GEN_3150;
  wire [31:0] _GEN_3151;
  wire [31:0] _GEN_3152;
  wire [31:0] _GEN_3153;
  wire [31:0] _GEN_3154;
  wire [31:0] _GEN_3155;
  wire [31:0] _GEN_3156;
  wire [31:0] _GEN_3157;
  wire [31:0] _GEN_3158;
  wire [31:0] _GEN_3159;
  wire [31:0] _GEN_3160;
  wire [31:0] _GEN_3161;
  wire [31:0] _GEN_3162;
  wire [31:0] _GEN_3163;
  wire [31:0] _GEN_3164;
  wire [31:0] _GEN_3165;
  wire [31:0] _GEN_3166;
  wire [31:0] _GEN_3167;
  wire [31:0] _GEN_3168;
  wire [31:0] _GEN_3169;
  wire [31:0] _GEN_3170;
  wire [31:0] _GEN_3171;
  wire [31:0] _GEN_3172;
  wire [31:0] _GEN_3173;
  wire [31:0] _GEN_3174;
  wire [31:0] _GEN_3175;
  wire [31:0] _GEN_3176;
  wire [31:0] _GEN_3177;
  wire [31:0] _GEN_3178;
  wire [31:0] _GEN_3179;
  wire [31:0] _GEN_3180;
  wire [31:0] _GEN_3181;
  wire [31:0] _GEN_3182;
  wire [31:0] _GEN_3183;
  wire [31:0] _GEN_3184;
  wire [31:0] _GEN_3185;
  wire [31:0] _GEN_3186;
  wire [31:0] _GEN_3187;
  wire [31:0] _GEN_3188;
  wire [31:0] _GEN_3189;
  wire [31:0] _GEN_3190;
  wire [31:0] _GEN_3191;
  wire [31:0] _GEN_3192;
  wire [31:0] _GEN_3193;
  wire [31:0] _GEN_3194;
  wire [31:0] _GEN_3195;
  wire [31:0] _GEN_3196;
  wire [31:0] _GEN_3197;
  wire [31:0] _GEN_3198;
  wire [31:0] _GEN_3199;
  wire [31:0] _GEN_3200;
  wire [31:0] _GEN_3201;
  wire [31:0] _GEN_3202;
  wire [31:0] _GEN_3203;
  wire [31:0] _GEN_3204;
  wire [31:0] _T_28888;
  wire [9:0] _T_28889;
  wire [1:0] _T_28890;
  wire [1:0] _T_28893_size;
  wire [9:0] _T_28893_source;
  RVX_MODULE_068 i_rvx_instance_31 (
    .rvx_port_2(rvx_signal_108),
    .rvx_port_0(rvx_signal_006),
    .rvx_port_4(rvx_signal_123),
    .rvx_port_5(rvx_signal_259),
    .rvx_port_1(rvx_signal_256),
    .rvx_port_3(rvx_signal_130)
  );
  RVX_MODULE_068 i_rvx_instance_29 (
    .rvx_port_2(rvx_signal_098),
    .rvx_port_0(rvx_signal_081),
    .rvx_port_4(rvx_signal_149),
    .rvx_port_5(rvx_signal_307),
    .rvx_port_1(rvx_signal_075),
    .rvx_port_3(rvx_signal_027)
  );
  RVX_MODULE_068 i_rvx_instance_02 (
    .rvx_port_2(rvx_signal_012),
    .rvx_port_0(rvx_signal_327),
    .rvx_port_4(rvx_signal_441),
    .rvx_port_5(rvx_signal_146),
    .rvx_port_1(rvx_signal_452),
    .rvx_port_3(rvx_signal_428)
  );
  RVX_MODULE_068 i_rvx_instance_27 (
    .rvx_port_2(rvx_signal_338),
    .rvx_port_0(rvx_signal_203),
    .rvx_port_4(rvx_signal_461),
    .rvx_port_5(rvx_signal_152),
    .rvx_port_1(rvx_signal_101),
    .rvx_port_3(rvx_signal_244)
  );
  RVX_MODULE_068 i_rvx_instance_23 (
    .rvx_port_2(rvx_signal_159),
    .rvx_port_0(rvx_signal_054),
    .rvx_port_4(rvx_signal_000),
    .rvx_port_5(rvx_signal_321),
    .rvx_port_1(rvx_signal_024),
    .rvx_port_3(rvx_signal_174)
  );
  RVX_MODULE_068 i_rvx_instance_15 (
    .rvx_port_2(rvx_signal_360),
    .rvx_port_0(rvx_signal_297),
    .rvx_port_4(rvx_signal_036),
    .rvx_port_5(rvx_signal_100),
    .rvx_port_1(rvx_signal_341),
    .rvx_port_3(rvx_signal_209)
  );
  RVX_MODULE_068 i_rvx_instance_07 (
    .rvx_port_2(rvx_signal_401),
    .rvx_port_0(rvx_signal_425),
    .rvx_port_4(rvx_signal_198),
    .rvx_port_5(rvx_signal_285),
    .rvx_port_1(rvx_signal_326),
    .rvx_port_3(rvx_signal_201)
  );
  RVX_MODULE_068 i_rvx_instance_26 (
    .rvx_port_2(rvx_signal_451),
    .rvx_port_0(rvx_signal_074),
    .rvx_port_4(rvx_signal_063),
    .rvx_port_5(rvx_signal_087),
    .rvx_port_1(rvx_signal_186),
    .rvx_port_3(rvx_signal_379)
  );
  RVX_MODULE_068 i_rvx_instance_32 (
    .rvx_port_2(rvx_signal_204),
    .rvx_port_0(rvx_signal_405),
    .rvx_port_4(rvx_signal_192),
    .rvx_port_5(rvx_signal_366),
    .rvx_port_1(rvx_signal_312),
    .rvx_port_3(rvx_signal_282)
  );
  RVX_MODULE_068 i_rvx_instance_18 (
    .rvx_port_2(rvx_signal_125),
    .rvx_port_0(rvx_signal_330),
    .rvx_port_4(rvx_signal_148),
    .rvx_port_5(rvx_signal_195),
    .rvx_port_1(rvx_signal_180),
    .rvx_port_3(rvx_signal_295)
  );
  RVX_MODULE_068 i_rvx_instance_14 (
    .rvx_port_2(rvx_signal_085),
    .rvx_port_0(rvx_signal_163),
    .rvx_port_4(rvx_signal_336),
    .rvx_port_5(rvx_signal_449),
    .rvx_port_1(rvx_signal_254),
    .rvx_port_3(rvx_signal_391)
  );
  RVX_MODULE_068 i_rvx_instance_21 (
    .rvx_port_2(rvx_signal_390),
    .rvx_port_0(rvx_signal_439),
    .rvx_port_4(rvx_signal_028),
    .rvx_port_5(rvx_signal_363),
    .rvx_port_1(rvx_signal_062),
    .rvx_port_3(rvx_signal_220)
  );
  RVX_MODULE_068 i_rvx_instance_22 (
    .rvx_port_2(rvx_signal_299),
    .rvx_port_0(rvx_signal_128),
    .rvx_port_4(rvx_signal_141),
    .rvx_port_5(rvx_signal_143),
    .rvx_port_1(rvx_signal_226),
    .rvx_port_3(rvx_signal_347)
  );
  RVX_MODULE_068 i_rvx_instance_25 (
    .rvx_port_2(rvx_signal_070),
    .rvx_port_0(rvx_signal_039),
    .rvx_port_4(rvx_signal_213),
    .rvx_port_5(rvx_signal_056),
    .rvx_port_1(rvx_signal_090),
    .rvx_port_3(rvx_signal_151)
  );
  RVX_MODULE_068 i_rvx_instance_16 (
    .rvx_port_2(rvx_signal_042),
    .rvx_port_0(rvx_signal_464),
    .rvx_port_4(rvx_signal_135),
    .rvx_port_5(rvx_signal_083),
    .rvx_port_1(rvx_signal_127),
    .rvx_port_3(rvx_signal_206)
  );
  RVX_MODULE_068 i_rvx_instance_04 (
    .rvx_port_2(rvx_signal_235),
    .rvx_port_0(rvx_signal_156),
    .rvx_port_4(rvx_signal_010),
    .rvx_port_5(rvx_signal_314),
    .rvx_port_1(rvx_signal_053),
    .rvx_port_3(rvx_signal_252)
  );
  RVX_MODULE_068 i_rvx_instance_33 (
    .rvx_port_2(rvx_signal_044),
    .rvx_port_0(rvx_signal_398),
    .rvx_port_4(rvx_signal_227),
    .rvx_port_5(rvx_signal_283),
    .rvx_port_1(rvx_signal_373),
    .rvx_port_3(rvx_signal_041)
  );
  RVX_MODULE_068 i_rvx_instance_01 (
    .rvx_port_2(rvx_signal_308),
    .rvx_port_0(rvx_signal_463),
    .rvx_port_4(rvx_signal_368),
    .rvx_port_5(rvx_signal_345),
    .rvx_port_1(rvx_signal_037),
    .rvx_port_3(rvx_signal_356)
  );
  RVX_MODULE_068 i_rvx_instance_06 (
    .rvx_port_2(rvx_signal_187),
    .rvx_port_0(rvx_signal_317),
    .rvx_port_4(rvx_signal_236),
    .rvx_port_5(rvx_signal_292),
    .rvx_port_1(rvx_signal_093),
    .rvx_port_3(rvx_signal_471)
  );
  RVX_MODULE_068 i_rvx_instance_12 (
    .rvx_port_2(rvx_signal_413),
    .rvx_port_0(rvx_signal_013),
    .rvx_port_4(rvx_signal_301),
    .rvx_port_5(rvx_signal_136),
    .rvx_port_1(rvx_signal_177),
    .rvx_port_3(rvx_signal_324)
  );
  RVX_MODULE_068 i_rvx_instance_11 (
    .rvx_port_2(rvx_signal_474),
    .rvx_port_0(rvx_signal_107),
    .rvx_port_4(rvx_signal_343),
    .rvx_port_5(rvx_signal_328),
    .rvx_port_1(rvx_signal_389),
    .rvx_port_3(rvx_signal_337)
  );
  RVX_MODULE_068 i_rvx_instance_08 (
    .rvx_port_2(rvx_signal_015),
    .rvx_port_0(rvx_signal_095),
    .rvx_port_4(rvx_signal_477),
    .rvx_port_5(rvx_signal_188),
    .rvx_port_1(rvx_signal_030),
    .rvx_port_3(rvx_signal_459)
  );
  RVX_MODULE_068 i_rvx_instance_09 (
    .rvx_port_2(rvx_signal_468),
    .rvx_port_0(rvx_signal_084),
    .rvx_port_4(rvx_signal_194),
    .rvx_port_5(rvx_signal_132),
    .rvx_port_1(rvx_signal_424),
    .rvx_port_3(rvx_signal_329)
  );
  RVX_MODULE_068 i_rvx_instance_03 (
    .rvx_port_2(rvx_signal_291),
    .rvx_port_0(rvx_signal_051),
    .rvx_port_4(rvx_signal_175),
    .rvx_port_5(rvx_signal_406),
    .rvx_port_1(rvx_signal_223),
    .rvx_port_3(rvx_signal_205)
  );
  RVX_MODULE_068 i_rvx_instance_30 (
    .rvx_port_2(rvx_signal_257),
    .rvx_port_0(rvx_signal_361),
    .rvx_port_4(rvx_signal_352),
    .rvx_port_5(rvx_signal_466),
    .rvx_port_1(rvx_signal_442),
    .rvx_port_3(rvx_signal_335)
  );
  RVX_MODULE_068 i_rvx_instance_24 (
    .rvx_port_2(rvx_signal_417),
    .rvx_port_0(rvx_signal_217),
    .rvx_port_4(rvx_signal_438),
    .rvx_port_5(rvx_signal_014),
    .rvx_port_1(rvx_signal_104),
    .rvx_port_3(rvx_signal_219)
  );
  RVX_MODULE_068 i_rvx_instance_20 (
    .rvx_port_2(rvx_signal_133),
    .rvx_port_0(rvx_signal_142),
    .rvx_port_4(rvx_signal_380),
    .rvx_port_5(rvx_signal_344),
    .rvx_port_1(rvx_signal_113),
    .rvx_port_3(rvx_signal_310)
  );
  RVX_MODULE_068 i_rvx_instance_17 (
    .rvx_port_2(rvx_signal_079),
    .rvx_port_0(rvx_signal_049),
    .rvx_port_4(rvx_signal_091),
    .rvx_port_5(rvx_signal_208),
    .rvx_port_1(rvx_signal_346),
    .rvx_port_3(rvx_signal_246)
  );
  RVX_MODULE_068 i_rvx_instance_10 (
    .rvx_port_2(rvx_signal_214),
    .rvx_port_0(rvx_signal_261),
    .rvx_port_4(rvx_signal_355),
    .rvx_port_5(rvx_signal_278),
    .rvx_port_1(rvx_signal_440),
    .rvx_port_3(rvx_signal_157)
  );
  RVX_MODULE_068 i_rvx_instance_13 (
    .rvx_port_2(rvx_signal_434),
    .rvx_port_0(rvx_signal_293),
    .rvx_port_4(rvx_signal_021),
    .rvx_port_5(rvx_signal_268),
    .rvx_port_1(rvx_signal_320),
    .rvx_port_3(rvx_signal_076)
  );
  RVX_MODULE_068 i_rvx_instance_28 (
    .rvx_port_2(rvx_signal_016),
    .rvx_port_0(rvx_signal_281),
    .rvx_port_4(rvx_signal_393),
    .rvx_port_5(rvx_signal_168),
    .rvx_port_1(rvx_signal_270),
    .rvx_port_3(rvx_signal_376)
  );
  RVX_MODULE_068 i_rvx_instance_19 (
    .rvx_port_2(rvx_signal_375),
    .rvx_port_0(rvx_signal_362),
    .rvx_port_4(rvx_signal_121),
    .rvx_port_5(rvx_signal_196),
    .rvx_port_1(rvx_signal_009),
    .rvx_port_3(rvx_signal_237)
  );
  RVX_MODULE_068 i_rvx_instance_05 (
    .rvx_port_2(rvx_signal_385),
    .rvx_port_0(rvx_signal_331),
    .rvx_port_4(rvx_signal_210),
    .rvx_port_5(rvx_signal_271),
    .rvx_port_1(rvx_signal_284),
    .rvx_port_3(rvx_signal_073)
  );
  RVX_MODULE_005 i_rvx_instance_00 (
    .rvx_port_05(rvx_signal_043),
    .rvx_port_15(rvx_signal_242),
    .rvx_port_04(rvx_signal_296),
    .rvx_port_03(rvx_signal_007),
    .rvx_port_07(rvx_signal_255),
    .rvx_port_06(rvx_signal_364),
    .rvx_port_14(rvx_signal_129),
    .rvx_port_12(rvx_signal_045),
    .rvx_port_13(rvx_signal_240),
    .rvx_port_00(rvx_signal_426),
    .rvx_port_01(rvx_signal_309),
    .rvx_port_08(rvx_signal_388),
    .rvx_port_11(rvx_signal_060),
    .rvx_port_02(rvx_signal_162),
    .rvx_port_10(rvx_signal_429),
    .rvx_port_09(rvx_signal_263)
  );
  assign _T_1259 = rvx_signal_065 & rvx_signal_099;
  assign _T_1260 = {_T_1259,rvx_signal_243};
  assign _T_1261 = rvx_signal_437 & rvx_signal_369;
  assign _T_1262 = {_T_1261,rvx_signal_057};
  assign _T_1263 = rvx_signal_382 & rvx_signal_221;
  assign _T_1264 = {_T_1263,rvx_signal_311};
  assign _T_1265 = rvx_signal_316 & rvx_signal_224;
  assign _T_1266 = {_T_1265,rvx_signal_089};
  assign _T_1267 = rvx_signal_165 & rvx_signal_066;
  assign _T_1268 = {_T_1267,rvx_signal_117};
  assign _T_1269 = rvx_signal_004 & rvx_signal_111;
  assign _T_1270 = {_T_1269,rvx_signal_116};
  assign _T_1271 = rvx_signal_272 & rvx_signal_179;
  assign _T_1272 = {_T_1271,rvx_signal_415};
  assign _T_1273 = rvx_signal_409 & rvx_signal_050;
  assign _T_1274 = {_T_1273,rvx_signal_289};
  assign _T_1275 = rvx_signal_202 & rvx_signal_215;
  assign _T_1276 = {_T_1275,rvx_signal_002};
  assign _T_1277 = rvx_signal_454 & rvx_signal_386;
  assign _T_1278 = {_T_1277,rvx_signal_395};
  assign _T_1279 = rvx_signal_092 & rvx_signal_450;
  assign _T_1280 = {_T_1279,rvx_signal_140};
  assign _T_1281 = rvx_signal_298 & rvx_signal_399;
  assign _T_1282 = {_T_1281,rvx_signal_023};
  assign _T_1283 = rvx_signal_096 & rvx_signal_067;
  assign _T_1284 = {_T_1283,rvx_signal_145};
  assign _T_1285 = rvx_signal_167 & rvx_signal_350;
  assign _T_1286 = {_T_1285,rvx_signal_025};
  assign _T_1287 = rvx_signal_294 & rvx_signal_265;
  assign _T_1288 = {_T_1287,rvx_signal_418};
  assign _T_1289 = rvx_signal_371 & rvx_signal_304;
  assign _T_1290 = {_T_1289,rvx_signal_008};
  assign _T_1291 = rvx_signal_103 & rvx_signal_058;
  assign _T_1292 = {_T_1291,rvx_signal_245};
  assign _T_1293 = rvx_signal_019 & rvx_signal_433;
  assign _T_1294 = {_T_1293,rvx_signal_114};
  assign _T_1295 = rvx_signal_080 & rvx_signal_465;
  assign _T_1296 = {_T_1295,rvx_signal_172};
  assign _T_1297 = rvx_signal_239 & rvx_signal_197;
  assign _T_1298 = {_T_1297,rvx_signal_266};
  assign _T_1299 = rvx_signal_124 & rvx_signal_358;
  assign _T_1300 = {_T_1299,rvx_signal_444};
  assign _T_1301 = rvx_signal_222 & rvx_signal_436;
  assign _T_1302 = {_T_1301,rvx_signal_088};
  assign _T_1303 = rvx_signal_306 & rvx_signal_001;
  assign _T_1304 = {_T_1303,rvx_signal_234};
  assign _T_1305 = rvx_signal_238 & rvx_signal_131;
  assign _T_1306 = {_T_1305,rvx_signal_097};
  assign _T_1307 = rvx_signal_011 & rvx_signal_410;
  assign _T_1308 = {_T_1307,rvx_signal_267};
  assign _T_1309 = rvx_signal_029 & rvx_signal_137;
  assign _T_1310 = {_T_1309,rvx_signal_248};
  assign _T_1311 = rvx_signal_166 & rvx_signal_178;
  assign _T_1312 = {_T_1311,rvx_signal_400};
  assign _T_1313 = rvx_signal_228 & rvx_signal_052;
  assign _T_1314 = {_T_1313,rvx_signal_430};
  assign _T_1315 = rvx_signal_183 & rvx_signal_423;
  assign _T_1316 = {_T_1315,rvx_signal_359};
  assign _T_1317 = rvx_signal_253 & rvx_signal_462;
  assign _T_1318 = {_T_1317,rvx_signal_332};
  assign _T_1319 = rvx_signal_033 & rvx_signal_475;
  assign _T_1320 = {_T_1319,rvx_signal_300};
  assign _T_1321 = rvx_signal_229 & rvx_signal_408;
  assign _T_1322 = {_T_1321,rvx_signal_032};
  assign _T_1325 = 4'h8 >= _T_1260;
  assign _T_1328 = _T_1325 ? 4'h8 : _T_1260;
  assign _T_1329 = _T_1325 ? 1'h0 : 1'h1;
  assign _T_1332 = _T_1262 >= _T_1264;
  assign _T_1335 = _T_1332 ? _T_1262 : _T_1264;
  assign _T_1336 = _T_1332 ? 1'h0 : 1'h1;
  assign _T_1337 = _T_1328 >= _T_1335;
  assign _GEN_3205 = {{1'd0}, _T_1336};
  assign _T_1339 = 2'h2 | _GEN_3205;
  assign _T_1340 = _T_1337 ? _T_1328 : _T_1335;
  assign _T_1341 = _T_1337 ? {{1'd0}, _T_1329} : _T_1339;
  assign _T_1344 = _T_1266 >= _T_1268;
  assign _T_1347 = _T_1344 ? _T_1266 : _T_1268;
  assign _T_1348 = _T_1344 ? 1'h0 : 1'h1;
  assign _T_1351 = _T_1270 >= _T_1272;
  assign _T_1354 = _T_1351 ? _T_1270 : _T_1272;
  assign _T_1355 = _T_1351 ? 1'h0 : 1'h1;
  assign _T_1356 = _T_1347 >= _T_1354;
  assign _GEN_3206 = {{1'd0}, _T_1355};
  assign _T_1358 = 2'h2 | _GEN_3206;
  assign _T_1359 = _T_1356 ? _T_1347 : _T_1354;
  assign _T_1360 = _T_1356 ? {{1'd0}, _T_1348} : _T_1358;
  assign _T_1361 = _T_1340 >= _T_1359;
  assign _GEN_3207 = {{1'd0}, _T_1360};
  assign _T_1363 = 3'h4 | _GEN_3207;
  assign _T_1364 = _T_1361 ? _T_1340 : _T_1359;
  assign _T_1365 = _T_1361 ? {{1'd0}, _T_1341} : _T_1363;
  assign _T_1368 = _T_1274 >= _T_1276;
  assign _T_1371 = _T_1368 ? _T_1274 : _T_1276;
  assign _T_1372 = _T_1368 ? 1'h0 : 1'h1;
  assign _T_1375 = _T_1278 >= _T_1280;
  assign _T_1378 = _T_1375 ? _T_1278 : _T_1280;
  assign _T_1379 = _T_1375 ? 1'h0 : 1'h1;
  assign _T_1380 = _T_1371 >= _T_1378;
  assign _GEN_3208 = {{1'd0}, _T_1379};
  assign _T_1382 = 2'h2 | _GEN_3208;
  assign _T_1383 = _T_1380 ? _T_1371 : _T_1378;
  assign _T_1384 = _T_1380 ? {{1'd0}, _T_1372} : _T_1382;
  assign _T_1387 = _T_1282 >= _T_1284;
  assign _T_1390 = _T_1387 ? _T_1282 : _T_1284;
  assign _T_1391 = _T_1387 ? 1'h0 : 1'h1;
  assign _T_1394 = _T_1286 >= _T_1288;
  assign _T_1397 = _T_1394 ? _T_1286 : _T_1288;
  assign _T_1398 = _T_1394 ? 1'h0 : 1'h1;
  assign _T_1399 = _T_1390 >= _T_1397;
  assign _GEN_3209 = {{1'd0}, _T_1398};
  assign _T_1401 = 2'h2 | _GEN_3209;
  assign _T_1402 = _T_1399 ? _T_1390 : _T_1397;
  assign _T_1403 = _T_1399 ? {{1'd0}, _T_1391} : _T_1401;
  assign _T_1404 = _T_1383 >= _T_1402;
  assign _GEN_3210 = {{1'd0}, _T_1403};
  assign _T_1406 = 3'h4 | _GEN_3210;
  assign _T_1407 = _T_1404 ? _T_1383 : _T_1402;
  assign _T_1408 = _T_1404 ? {{1'd0}, _T_1384} : _T_1406;
  assign _T_1409 = _T_1364 >= _T_1407;
  assign _GEN_3211 = {{1'd0}, _T_1408};
  assign _T_1411 = 4'h8 | _GEN_3211;
  assign _T_1412 = _T_1409 ? _T_1364 : _T_1407;
  assign _T_1413 = _T_1409 ? {{1'd0}, _T_1365} : _T_1411;
  assign _T_1416 = _T_1290 >= _T_1292;
  assign _T_1419 = _T_1416 ? _T_1290 : _T_1292;
  assign _T_1420 = _T_1416 ? 1'h0 : 1'h1;
  assign _T_1423 = _T_1294 >= _T_1296;
  assign _T_1426 = _T_1423 ? _T_1294 : _T_1296;
  assign _T_1427 = _T_1423 ? 1'h0 : 1'h1;
  assign _T_1428 = _T_1419 >= _T_1426;
  assign _GEN_3212 = {{1'd0}, _T_1427};
  assign _T_1430 = 2'h2 | _GEN_3212;
  assign _T_1431 = _T_1428 ? _T_1419 : _T_1426;
  assign _T_1432 = _T_1428 ? {{1'd0}, _T_1420} : _T_1430;
  assign _T_1435 = _T_1298 >= _T_1300;
  assign _T_1438 = _T_1435 ? _T_1298 : _T_1300;
  assign _T_1439 = _T_1435 ? 1'h0 : 1'h1;
  assign _T_1442 = _T_1302 >= _T_1304;
  assign _T_1445 = _T_1442 ? _T_1302 : _T_1304;
  assign _T_1446 = _T_1442 ? 1'h0 : 1'h1;
  assign _T_1447 = _T_1438 >= _T_1445;
  assign _GEN_3213 = {{1'd0}, _T_1446};
  assign _T_1449 = 2'h2 | _GEN_3213;
  assign _T_1450 = _T_1447 ? _T_1438 : _T_1445;
  assign _T_1451 = _T_1447 ? {{1'd0}, _T_1439} : _T_1449;
  assign _T_1452 = _T_1431 >= _T_1450;
  assign _GEN_3214 = {{1'd0}, _T_1451};
  assign _T_1454 = 3'h4 | _GEN_3214;
  assign _T_1455 = _T_1452 ? _T_1431 : _T_1450;
  assign _T_1456 = _T_1452 ? {{1'd0}, _T_1432} : _T_1454;
  assign _T_1459 = _T_1306 >= _T_1308;
  assign _T_1462 = _T_1459 ? _T_1306 : _T_1308;
  assign _T_1463 = _T_1459 ? 1'h0 : 1'h1;
  assign _T_1466 = _T_1310 >= _T_1312;
  assign _T_1469 = _T_1466 ? _T_1310 : _T_1312;
  assign _T_1470 = _T_1466 ? 1'h0 : 1'h1;
  assign _T_1471 = _T_1462 >= _T_1469;
  assign _GEN_3215 = {{1'd0}, _T_1470};
  assign _T_1473 = 2'h2 | _GEN_3215;
  assign _T_1474 = _T_1471 ? _T_1462 : _T_1469;
  assign _T_1475 = _T_1471 ? {{1'd0}, _T_1463} : _T_1473;
  assign _T_1478 = _T_1314 >= _T_1316;
  assign _T_1481 = _T_1478 ? _T_1314 : _T_1316;
  assign _T_1482 = _T_1478 ? 1'h0 : 1'h1;
  assign _T_1485 = _T_1318 >= _T_1320;
  assign _T_1488 = _T_1485 ? _T_1318 : _T_1320;
  assign _T_1489 = _T_1485 ? 1'h0 : 1'h1;
  assign _T_1490 = _T_1481 >= _T_1488;
  assign _GEN_3216 = {{1'd0}, _T_1489};
  assign _T_1492 = 2'h2 | _GEN_3216;
  assign _T_1493 = _T_1490 ? _T_1481 : _T_1488;
  assign _T_1494 = _T_1490 ? {{1'd0}, _T_1482} : _T_1492;
  assign _T_1495 = _T_1474 >= _T_1493;
  assign _GEN_3217 = {{1'd0}, _T_1494};
  assign _T_1497 = 3'h4 | _GEN_3217;
  assign _T_1498 = _T_1495 ? _T_1474 : _T_1493;
  assign _T_1499 = _T_1495 ? {{1'd0}, _T_1475} : _T_1497;
  assign _T_1500 = _T_1455 >= _T_1498;
  assign _GEN_3218 = {{1'd0}, _T_1499};
  assign _T_1502 = 4'h8 | _GEN_3218;
  assign _T_1503 = _T_1500 ? _T_1455 : _T_1498;
  assign _T_1504 = _T_1500 ? {{1'd0}, _T_1456} : _T_1502;
  assign _T_1505 = _T_1412 >= _T_1503;
  assign _GEN_3219 = {{1'd0}, _T_1504};
  assign _T_1507 = 5'h10 | _GEN_3219;
  assign _T_1508 = _T_1505 ? _T_1412 : _T_1503;
  assign _T_1509 = _T_1505 ? {{1'd0}, _T_1413} : _T_1507;
  assign _T_1511 = _T_1508 >= _T_1322;
  assign _T_1514 = _T_1511 ? _T_1508 : _T_1322;
  assign _T_1515 = _T_1511 ? {{1'd0}, _T_1509} : 6'h20;
  assign _T_1519 = {1'h1,rvx_signal_435};
  assign _T_1520 = _T_1517 > _T_1519;
  assign _T_1529 = rvx_signal_189 - 1'h1;
  assign _T_1530 = $unsigned(_T_1529);
  assign _T_1531 = _T_1530[0:0];
  assign _T_1532 = rvx_signal_189 & _T_1531;
  assign _T_1534 = _T_1532 == 1'h0;
  assign _T_1536 = _T_1534 | rvx_port_41;
  assign _T_1538 = _T_1536 == 1'h0;
  assign _T_1541 = 64'h1 << rvx_signal_153;
  assign _T_1542 = _T_1541[32:0];
  assign _T_1544 = rvx_signal_189 ? _T_1542 : 33'h0;
  assign _T_1551 = rvx_signal_161[1];
  assign _T_1552 = rvx_signal_161[2];
  assign _T_1553 = rvx_signal_161[3];
  assign _T_1554 = rvx_signal_161[4];
  assign _T_1555 = rvx_signal_161[5];
  assign _T_1556 = rvx_signal_161[6];
  assign _T_1557 = rvx_signal_161[7];
  assign _T_1558 = rvx_signal_161[8];
  assign _T_1559 = rvx_signal_161[9];
  assign _T_1560 = rvx_signal_161[10];
  assign _T_1561 = rvx_signal_161[11];
  assign _T_1562 = rvx_signal_161[12];
  assign _T_1563 = rvx_signal_161[13];
  assign _T_1564 = rvx_signal_161[14];
  assign _T_1565 = rvx_signal_161[15];
  assign _T_1566 = rvx_signal_161[16];
  assign _T_1567 = rvx_signal_161[17];
  assign _T_1568 = rvx_signal_161[18];
  assign _T_1569 = rvx_signal_161[19];
  assign _T_1570 = rvx_signal_161[20];
  assign _T_1571 = rvx_signal_161[21];
  assign _T_1572 = rvx_signal_161[22];
  assign _T_1573 = rvx_signal_161[23];
  assign _T_1574 = rvx_signal_161[24];
  assign _T_1575 = rvx_signal_161[25];
  assign _T_1576 = rvx_signal_161[26];
  assign _T_1577 = rvx_signal_161[27];
  assign _T_1578 = rvx_signal_161[28];
  assign _T_1579 = rvx_signal_161[29];
  assign _T_1580 = rvx_signal_161[30];
  assign _T_1581 = rvx_signal_161[31];
  assign _T_1582 = rvx_signal_161[32];
  assign _T_1626 = rvx_signal_065 == 1'h0;
  assign _T_1627 = rvx_signal_017 | rvx_signal_269;
  assign _T_1629 = rvx_signal_017 == 1'h0;
  assign _GEN_8 = _T_1627 ? _T_1629 : rvx_signal_065;
  assign _T_1631 = rvx_signal_437 == 1'h0;
  assign _T_1632 = rvx_signal_164 | rvx_signal_119;
  assign _T_1634 = rvx_signal_164 == 1'h0;
  assign _GEN_9 = _T_1632 ? _T_1634 : rvx_signal_437;
  assign _T_1636 = rvx_signal_382 == 1'h0;
  assign _T_1637 = rvx_signal_427 | rvx_signal_184;
  assign _T_1639 = rvx_signal_427 == 1'h0;
  assign _GEN_10 = _T_1637 ? _T_1639 : rvx_signal_382;
  assign _T_1641 = rvx_signal_316 == 1'h0;
  assign _T_1642 = rvx_signal_005 | rvx_signal_251;
  assign _T_1644 = rvx_signal_005 == 1'h0;
  assign _GEN_11 = _T_1642 ? _T_1644 : rvx_signal_316;
  assign _T_1646 = rvx_signal_165 == 1'h0;
  assign _T_1647 = rvx_signal_275 | rvx_signal_199;
  assign _T_1649 = rvx_signal_275 == 1'h0;
  assign _GEN_12 = _T_1647 ? _T_1649 : rvx_signal_165;
  assign _T_1651 = rvx_signal_004 == 1'h0;
  assign _T_1652 = rvx_signal_182 | rvx_signal_378;
  assign _T_1654 = rvx_signal_182 == 1'h0;
  assign _GEN_13 = _T_1652 ? _T_1654 : rvx_signal_004;
  assign _T_1656 = rvx_signal_272 == 1'h0;
  assign _T_1657 = rvx_signal_185 | rvx_signal_349;
  assign _T_1659 = rvx_signal_185 == 1'h0;
  assign _GEN_14 = _T_1657 ? _T_1659 : rvx_signal_272;
  assign _T_1661 = rvx_signal_409 == 1'h0;
  assign _T_1662 = rvx_signal_110 | rvx_signal_241;
  assign _T_1664 = rvx_signal_110 == 1'h0;
  assign _GEN_15 = _T_1662 ? _T_1664 : rvx_signal_409;
  assign _T_1666 = rvx_signal_202 == 1'h0;
  assign _T_1667 = rvx_signal_372 | rvx_signal_365;
  assign _T_1669 = rvx_signal_372 == 1'h0;
  assign _GEN_16 = _T_1667 ? _T_1669 : rvx_signal_202;
  assign _T_1671 = rvx_signal_454 == 1'h0;
  assign _T_1672 = rvx_signal_290 | rvx_signal_422;
  assign _T_1674 = rvx_signal_290 == 1'h0;
  assign _GEN_17 = _T_1672 ? _T_1674 : rvx_signal_454;
  assign _T_1676 = rvx_signal_092 == 1'h0;
  assign _T_1677 = rvx_signal_407 | rvx_signal_351;
  assign _T_1679 = rvx_signal_407 == 1'h0;
  assign _GEN_18 = _T_1677 ? _T_1679 : rvx_signal_092;
  assign _T_1681 = rvx_signal_298 == 1'h0;
  assign _T_1682 = rvx_signal_126 | rvx_signal_068;
  assign _T_1684 = rvx_signal_126 == 1'h0;
  assign _GEN_19 = _T_1682 ? _T_1684 : rvx_signal_298;
  assign _T_1686 = rvx_signal_096 == 1'h0;
  assign _T_1687 = rvx_signal_374 | rvx_signal_118;
  assign _T_1689 = rvx_signal_374 == 1'h0;
  assign _GEN_20 = _T_1687 ? _T_1689 : rvx_signal_096;
  assign _T_1691 = rvx_signal_167 == 1'h0;
  assign _T_1692 = rvx_signal_318 | rvx_signal_305;
  assign _T_1694 = rvx_signal_318 == 1'h0;
  assign _GEN_21 = _T_1692 ? _T_1694 : rvx_signal_167;
  assign _T_1696 = rvx_signal_294 == 1'h0;
  assign _T_1697 = rvx_signal_279 | rvx_signal_233;
  assign _T_1699 = rvx_signal_279 == 1'h0;
  assign _GEN_22 = _T_1697 ? _T_1699 : rvx_signal_294;
  assign _T_1701 = rvx_signal_371 == 1'h0;
  assign _T_1702 = rvx_signal_303 | rvx_signal_022;
  assign _T_1704 = rvx_signal_303 == 1'h0;
  assign _GEN_23 = _T_1702 ? _T_1704 : rvx_signal_371;
  assign _T_1706 = rvx_signal_103 == 1'h0;
  assign _T_1707 = rvx_signal_038 | rvx_signal_086;
  assign _T_1709 = rvx_signal_038 == 1'h0;
  assign _GEN_24 = _T_1707 ? _T_1709 : rvx_signal_103;
  assign _T_1711 = rvx_signal_019 == 1'h0;
  assign _T_1712 = rvx_signal_077 | rvx_signal_416;
  assign _T_1714 = rvx_signal_077 == 1'h0;
  assign _GEN_25 = _T_1712 ? _T_1714 : rvx_signal_019;
  assign _T_1716 = rvx_signal_080 == 1'h0;
  assign _T_1717 = rvx_signal_384 | rvx_signal_190;
  assign _T_1719 = rvx_signal_384 == 1'h0;
  assign _GEN_26 = _T_1717 ? _T_1719 : rvx_signal_080;
  assign _T_1721 = rvx_signal_239 == 1'h0;
  assign _T_1722 = rvx_signal_446 | rvx_signal_225;
  assign _T_1724 = rvx_signal_446 == 1'h0;
  assign _GEN_27 = _T_1722 ? _T_1724 : rvx_signal_239;
  assign _T_1726 = rvx_signal_124 == 1'h0;
  assign _T_1727 = rvx_signal_443 | rvx_signal_469;
  assign _T_1729 = rvx_signal_443 == 1'h0;
  assign _GEN_28 = _T_1727 ? _T_1729 : rvx_signal_124;
  assign _T_1731 = rvx_signal_222 == 1'h0;
  assign _T_1732 = rvx_signal_150 | rvx_signal_460;
  assign _T_1734 = rvx_signal_150 == 1'h0;
  assign _GEN_29 = _T_1732 ? _T_1734 : rvx_signal_222;
  assign _T_1736 = rvx_signal_306 == 1'h0;
  assign _T_1737 = rvx_signal_383 | rvx_signal_404;
  assign _T_1739 = rvx_signal_383 == 1'h0;
  assign _GEN_30 = _T_1737 ? _T_1739 : rvx_signal_306;
  assign _T_1741 = rvx_signal_238 == 1'h0;
  assign _T_1742 = rvx_signal_048 | rvx_signal_315;
  assign _T_1744 = rvx_signal_048 == 1'h0;
  assign _GEN_31 = _T_1742 ? _T_1744 : rvx_signal_238;
  assign _T_1746 = rvx_signal_011 == 1'h0;
  assign _T_1747 = rvx_signal_249 | rvx_signal_003;
  assign _T_1749 = rvx_signal_249 == 1'h0;
  assign _GEN_32 = _T_1747 ? _T_1749 : rvx_signal_011;
  assign _T_1751 = rvx_signal_029 == 1'h0;
  assign _T_1752 = rvx_signal_064 | rvx_signal_181;
  assign _T_1754 = rvx_signal_064 == 1'h0;
  assign _GEN_33 = _T_1752 ? _T_1754 : rvx_signal_029;
  assign _T_1756 = rvx_signal_166 == 1'h0;
  assign _T_1757 = rvx_signal_470 | rvx_signal_287;
  assign _T_1759 = rvx_signal_470 == 1'h0;
  assign _GEN_34 = _T_1757 ? _T_1759 : rvx_signal_166;
  assign _T_1761 = rvx_signal_228 == 1'h0;
  assign _T_1762 = rvx_signal_258 | rvx_signal_072;
  assign _T_1764 = rvx_signal_258 == 1'h0;
  assign _GEN_35 = _T_1762 ? _T_1764 : rvx_signal_228;
  assign _T_1766 = rvx_signal_183 == 1'h0;
  assign _T_1767 = rvx_signal_034 | rvx_signal_276;
  assign _T_1769 = rvx_signal_034 == 1'h0;
  assign _GEN_36 = _T_1767 ? _T_1769 : rvx_signal_183;
  assign _T_1771 = rvx_signal_253 == 1'h0;
  assign _T_1772 = rvx_signal_018 | rvx_signal_273;
  assign _T_1774 = rvx_signal_018 == 1'h0;
  assign _GEN_37 = _T_1772 ? _T_1774 : rvx_signal_253;
  assign _T_1776 = rvx_signal_033 == 1'h0;
  assign _T_1777 = rvx_signal_155 | rvx_signal_445;
  assign _T_1779 = rvx_signal_155 == 1'h0;
  assign _GEN_38 = _T_1777 ? _T_1779 : rvx_signal_033;
  assign _T_1781 = rvx_signal_229 == 1'h0;
  assign _T_1782 = rvx_signal_144 | rvx_signal_173;
  assign _T_1784 = rvx_signal_144 == 1'h0;
  assign _GEN_39 = _T_1782 ? _T_1784 : rvx_signal_229;
  assign _T_1792 = rvx_signal_431 - 1'h1;
  assign _T_1793 = $unsigned(_T_1792);
  assign _T_1794 = _T_1793[0:0];
  assign _T_1795 = rvx_signal_431 & _T_1794;
  assign _T_1797 = _T_1795 == 1'h0;
  assign _T_1799 = _T_1797 | rvx_port_41;
  assign _T_1801 = _T_1799 == 1'h0;
  assign _T_1805 = 64'h1 << rvx_signal_120;
  assign _T_1806 = _T_1805[32:0];
  assign rvx_signal_432 = rvx_signal_431 ? _T_1806 : 33'h0;
  assign _T_1808 = rvx_signal_432[0];
  assign _T_1809 = rvx_signal_432[1];
  assign _T_1810 = rvx_signal_432[2];
  assign _T_1811 = rvx_signal_432[3];
  assign _T_1812 = rvx_signal_432[4];
  assign _T_1813 = rvx_signal_432[5];
  assign _T_1814 = rvx_signal_432[6];
  assign _T_1815 = rvx_signal_432[7];
  assign _T_1816 = rvx_signal_432[8];
  assign _T_1817 = rvx_signal_432[9];
  assign _T_1818 = rvx_signal_432[10];
  assign _T_1819 = rvx_signal_432[11];
  assign _T_1820 = rvx_signal_432[12];
  assign _T_1821 = rvx_signal_432[13];
  assign _T_1822 = rvx_signal_432[14];
  assign _T_1823 = rvx_signal_432[15];
  assign _T_1824 = rvx_signal_432[16];
  assign _T_1825 = rvx_signal_432[17];
  assign _T_1826 = rvx_signal_432[18];
  assign _T_1827 = rvx_signal_432[19];
  assign _T_1828 = rvx_signal_432[20];
  assign _T_1829 = rvx_signal_432[21];
  assign _T_1830 = rvx_signal_432[22];
  assign _T_1831 = rvx_signal_432[23];
  assign _T_1832 = rvx_signal_432[24];
  assign _T_1833 = rvx_signal_432[25];
  assign _T_1834 = rvx_signal_432[26];
  assign _T_1835 = rvx_signal_432[27];
  assign _T_1836 = rvx_signal_432[28];
  assign _T_1837 = rvx_signal_432[29];
  assign _T_1838 = rvx_signal_432[30];
  assign _T_1839 = rvx_signal_432[31];
  assign _T_1840 = rvx_signal_432[32];
  assign _T_1851 = _T_31_a_bits_opcode == 3'h4;
  assign _T_1852 = _T_31_a_bits_address[27:2];
  assign _T_1853 = {_T_31_a_bits_source,_T_31_a_bits_size};
  assign _T_2903 = rvx_signal_060 ^ 24'h400;
  assign _T_2904 = _T_2903 & 24'hf7f3c0;
  assign _T_2906 = _T_2904 == 24'h0;
  assign _T_2912 = rvx_signal_060;
  assign _T_2913 = _T_2912 & 24'hf7f3c0;
  assign _T_2915 = _T_2913 == 24'h0;
  assign _T_2921 = rvx_signal_060 ^ 24'h5;
  assign _T_2922 = _T_2921 & 24'hf7f3c0;
  assign _T_2924 = _T_2922 == 24'h0;
  assign _T_2930 = rvx_signal_060 ^ 24'ha;
  assign _T_2931 = _T_2930 & 24'hf7f3c0;
  assign _T_2933 = _T_2931 == 24'h0;
  assign _T_2939 = rvx_signal_060 ^ 24'h18;
  assign _T_2940 = _T_2939 & 24'hf7f3c0;
  assign _T_2942 = _T_2940 == 24'h0;
  assign _T_2948 = rvx_signal_060 ^ 24'h19;
  assign _T_2949 = _T_2948 & 24'hf7f3c0;
  assign _T_2951 = _T_2949 == 24'h0;
  assign _T_2957 = rvx_signal_060 ^ 24'he;
  assign _T_2958 = _T_2957 & 24'hf7f3c0;
  assign _T_2960 = _T_2958 == 24'h0;
  assign _T_2966 = rvx_signal_060 ^ 24'h14;
  assign _T_2967 = _T_2966 & 24'hf7f3c0;
  assign _T_2969 = _T_2967 == 24'h0;
  assign _T_2975 = rvx_signal_060 ^ 24'h801;
  assign _T_2976 = _T_2975 & 24'hf7f3c0;
  assign _T_2978 = _T_2976 == 24'h0;
  assign _T_2984 = rvx_signal_060 ^ 24'h1d;
  assign _T_2985 = _T_2984 & 24'hf7f3c0;
  assign _T_2987 = _T_2985 == 24'h0;
  assign _T_2993 = rvx_signal_060 ^ 24'h80001;
  assign _T_2994 = _T_2993 & 24'hf7f3c0;
  assign _T_2996 = _T_2994 == 24'h0;
  assign _T_3002 = rvx_signal_060 ^ 24'h1;
  assign _T_3003 = _T_3002 & 24'hf7f3c0;
  assign _T_3005 = _T_3003 == 24'h0;
  assign _T_3011 = rvx_signal_060 ^ 24'h6;
  assign _T_3012 = _T_3011 & 24'hf7f3c0;
  assign _T_3014 = _T_3012 == 24'h0;
  assign _T_3020 = rvx_signal_060 ^ 24'h1c;
  assign _T_3021 = _T_3020 & 24'hf7f3c0;
  assign _T_3023 = _T_3021 == 24'h0;
  assign _T_3029 = rvx_signal_060 ^ 24'h15;
  assign _T_3030 = _T_3029 & 24'hf7f3c0;
  assign _T_3032 = _T_3030 == 24'h0;
  assign _T_3038 = rvx_signal_060 ^ 24'h9;
  assign _T_3039 = _T_3038 & 24'hf7f3c0;
  assign _T_3041 = _T_3039 == 24'h0;
  assign _T_3047 = rvx_signal_060 ^ 24'hd;
  assign _T_3048 = _T_3047 & 24'hf7f3c0;
  assign _T_3050 = _T_3048 == 24'h0;
  assign _T_3056 = rvx_signal_060 ^ 24'h2;
  assign _T_3057 = _T_3056 & 24'hf7f3c0;
  assign _T_3059 = _T_3057 == 24'h0;
  assign _T_3065 = rvx_signal_060 ^ 24'h20;
  assign _T_3066 = _T_3065 & 24'hf7f3c0;
  assign _T_3068 = _T_3066 == 24'h0;
  assign _T_3074 = rvx_signal_060 ^ 24'h11;
  assign _T_3075 = _T_3074 & 24'hf7f3c0;
  assign _T_3077 = _T_3075 == 24'h0;
  assign _T_3083 = rvx_signal_060 ^ 24'h80000;
  assign _T_3084 = _T_3083 & 24'hf7f3c0;
  assign _T_3086 = _T_3084 == 24'h0;
  assign _T_3092 = rvx_signal_060 ^ 24'h800;
  assign _T_3093 = _T_3092 & 24'hf7f3c0;
  assign _T_3095 = _T_3093 == 24'h0;
  assign _T_3101 = rvx_signal_060 ^ 24'h16;
  assign _T_3102 = _T_3101 & 24'hf7f3c0;
  assign _T_3104 = _T_3102 == 24'h0;
  assign _T_3110 = rvx_signal_060 ^ 24'h1b;
  assign _T_3111 = _T_3110 & 24'hf7f3c0;
  assign _T_3113 = _T_3111 == 24'h0;
  assign _T_3119 = rvx_signal_060 ^ 24'hc;
  assign _T_3120 = _T_3119 & 24'hf7f3c0;
  assign _T_3122 = _T_3120 == 24'h0;
  assign _T_3128 = rvx_signal_060 ^ 24'h7;
  assign _T_3129 = _T_3128 & 24'hf7f3c0;
  assign _T_3131 = _T_3129 == 24'h0;
  assign _T_3137 = rvx_signal_060 ^ 24'h3;
  assign _T_3138 = _T_3137 & 24'hf7f3c0;
  assign _T_3140 = _T_3138 == 24'h0;
  assign _T_3146 = rvx_signal_060 ^ 24'h401;
  assign _T_3147 = _T_3146 & 24'hf7f3c0;
  assign _T_3149 = _T_3147 == 24'h0;
  assign _T_3155 = rvx_signal_060 ^ 24'h12;
  assign _T_3156 = _T_3155 & 24'hf7f3c0;
  assign _T_3158 = _T_3156 == 24'h0;
  assign _T_3164 = rvx_signal_060 ^ 24'h10;
  assign _T_3165 = _T_3164 & 24'hf7f3c0;
  assign _T_3167 = _T_3165 == 24'h0;
  assign _T_3173 = rvx_signal_060 ^ 24'h1f;
  assign _T_3174 = _T_3173 & 24'hf7f3c0;
  assign _T_3176 = _T_3174 == 24'h0;
  assign _T_3182 = rvx_signal_060 ^ 24'hb;
  assign _T_3183 = _T_3182 & 24'hf7f3c0;
  assign _T_3185 = _T_3183 == 24'h0;
  assign _T_3191 = rvx_signal_060 ^ 24'h1a;
  assign _T_3192 = _T_3191 & 24'hf7f3c0;
  assign _T_3194 = _T_3192 == 24'h0;
  assign _T_3200 = rvx_signal_060 ^ 24'h17;
  assign _T_3201 = _T_3200 & 24'hf7f3c0;
  assign _T_3203 = _T_3201 == 24'h0;
  assign _T_3209 = rvx_signal_060 ^ 24'h8;
  assign _T_3210 = _T_3209 & 24'hf7f3c0;
  assign _T_3212 = _T_3210 == 24'h0;
  assign _T_3218 = rvx_signal_060 ^ 24'h1e;
  assign _T_3219 = _T_3218 & 24'hf7f3c0;
  assign _T_3221 = _T_3219 == 24'h0;
  assign _T_3227 = rvx_signal_060 ^ 24'h13;
  assign _T_3228 = _T_3227 & 24'hf7f3c0;
  assign _T_3230 = _T_3228 == 24'h0;
  assign _T_3236 = rvx_signal_060 ^ 24'h4;
  assign _T_3237 = _T_3236 & 24'hf7f3c0;
  assign _T_3239 = _T_3237 == 24'h0;
  assign _T_3245 = rvx_signal_060 ^ 24'hf;
  assign _T_3246 = _T_3245 & 24'hf7f3c0;
  assign _T_3248 = _T_3246 == 24'h0;
  assign _T_4212 = rvx_signal_429[0];
  assign _T_4213 = rvx_signal_429[1];
  assign _T_4214 = rvx_signal_429[2];
  assign _T_4215 = rvx_signal_429[3];
  assign _T_4219 = _T_4212 ? 8'hff : 8'h0;
  assign _T_4223 = _T_4213 ? 8'hff : 8'h0;
  assign _T_4227 = _T_4214 ? 8'hff : 8'h0;
  assign _T_4231 = _T_4215 ? 8'hff : 8'h0;
  assign _T_4232 = {_T_4223,_T_4219};
  assign _T_4233 = {_T_4231,_T_4227};
  assign _T_4234 = {_T_4233,_T_4232};
  assign _T_4242 = _T_4234[0];
  assign _T_4246 = ~ _T_4242;
  assign _T_4248 = _T_4246 == 1'h0;
  assign _T_4255 = rvx_signal_162[0];
  assign _T_4282 = _T_4234[1];
  assign _T_4286 = ~ _T_4282;
  assign _T_4288 = _T_4286 == 1'h0;
  assign _T_4295 = rvx_signal_162[1];
  assign _GEN_3220 = {{1'd0}, rvx_signal_065};
  assign _T_4310 = _GEN_3220 << 1;
  assign _T_4322 = _T_4234[2];
  assign _T_4326 = ~ _T_4322;
  assign _T_4328 = _T_4326 == 1'h0;
  assign _T_4335 = rvx_signal_162[2];
  assign _GEN_3221 = {{2'd0}, rvx_signal_437};
  assign _T_4350 = _GEN_3221 << 2;
  assign _GEN_3222 = {{1'd0}, _T_4310};
  assign _T_4354 = _GEN_3222 | _T_4350;
  assign _T_4362 = _T_4234[3];
  assign _T_4366 = ~ _T_4362;
  assign _T_4368 = _T_4366 == 1'h0;
  assign _T_4375 = rvx_signal_162[3];
  assign _GEN_3223 = {{3'd0}, rvx_signal_382};
  assign _T_4390 = _GEN_3223 << 3;
  assign _GEN_3224 = {{1'd0}, _T_4354};
  assign _T_4394 = _GEN_3224 | _T_4390;
  assign _T_4402 = _T_4234[4];
  assign _T_4406 = ~ _T_4402;
  assign _T_4408 = _T_4406 == 1'h0;
  assign _T_4415 = rvx_signal_162[4];
  assign _GEN_3225 = {{4'd0}, rvx_signal_316};
  assign _T_4430 = _GEN_3225 << 4;
  assign _GEN_3226 = {{1'd0}, _T_4394};
  assign _T_4434 = _GEN_3226 | _T_4430;
  assign _T_4442 = _T_4234[5];
  assign _T_4446 = ~ _T_4442;
  assign _T_4448 = _T_4446 == 1'h0;
  assign _T_4455 = rvx_signal_162[5];
  assign _GEN_3227 = {{5'd0}, rvx_signal_165};
  assign _T_4470 = _GEN_3227 << 5;
  assign _GEN_3228 = {{1'd0}, _T_4434};
  assign _T_4474 = _GEN_3228 | _T_4470;
  assign _T_4482 = _T_4234[6];
  assign _T_4486 = ~ _T_4482;
  assign _T_4488 = _T_4486 == 1'h0;
  assign _T_4495 = rvx_signal_162[6];
  assign _GEN_3229 = {{6'd0}, rvx_signal_004};
  assign _T_4510 = _GEN_3229 << 6;
  assign _GEN_3230 = {{1'd0}, _T_4474};
  assign _T_4514 = _GEN_3230 | _T_4510;
  assign _T_4522 = _T_4234[7];
  assign _T_4526 = ~ _T_4522;
  assign _T_4528 = _T_4526 == 1'h0;
  assign _T_4535 = rvx_signal_162[7];
  assign _GEN_3231 = {{7'd0}, rvx_signal_272};
  assign _T_4550 = _GEN_3231 << 7;
  assign _GEN_3232 = {{1'd0}, _T_4514};
  assign _T_4554 = _GEN_3232 | _T_4550;
  assign _T_4562 = _T_4234[8];
  assign _T_4566 = ~ _T_4562;
  assign _T_4568 = _T_4566 == 1'h0;
  assign _T_4575 = rvx_signal_162[8];
  assign _GEN_3233 = {{8'd0}, rvx_signal_409};
  assign _T_4590 = _GEN_3233 << 8;
  assign _GEN_3234 = {{1'd0}, _T_4554};
  assign _T_4594 = _GEN_3234 | _T_4590;
  assign _T_4602 = _T_4234[9];
  assign _T_4606 = ~ _T_4602;
  assign _T_4608 = _T_4606 == 1'h0;
  assign _T_4615 = rvx_signal_162[9];
  assign _GEN_3235 = {{9'd0}, rvx_signal_202};
  assign _T_4630 = _GEN_3235 << 9;
  assign _GEN_3236 = {{1'd0}, _T_4594};
  assign _T_4634 = _GEN_3236 | _T_4630;
  assign _T_4642 = _T_4234[10];
  assign _T_4646 = ~ _T_4642;
  assign _T_4648 = _T_4646 == 1'h0;
  assign _T_4655 = rvx_signal_162[10];
  assign _GEN_3237 = {{10'd0}, rvx_signal_454};
  assign _T_4670 = _GEN_3237 << 10;
  assign _GEN_3238 = {{1'd0}, _T_4634};
  assign _T_4674 = _GEN_3238 | _T_4670;
  assign _T_4682 = _T_4234[11];
  assign _T_4686 = ~ _T_4682;
  assign _T_4688 = _T_4686 == 1'h0;
  assign _T_4695 = rvx_signal_162[11];
  assign _GEN_3239 = {{11'd0}, rvx_signal_092};
  assign _T_4710 = _GEN_3239 << 11;
  assign _GEN_3240 = {{1'd0}, _T_4674};
  assign _T_4714 = _GEN_3240 | _T_4710;
  assign _T_4722 = _T_4234[12];
  assign _T_4726 = ~ _T_4722;
  assign _T_4728 = _T_4726 == 1'h0;
  assign _T_4735 = rvx_signal_162[12];
  assign _GEN_3241 = {{12'd0}, rvx_signal_298};
  assign _T_4750 = _GEN_3241 << 12;
  assign _GEN_3242 = {{1'd0}, _T_4714};
  assign _T_4754 = _GEN_3242 | _T_4750;
  assign _T_4762 = _T_4234[13];
  assign _T_4766 = ~ _T_4762;
  assign _T_4768 = _T_4766 == 1'h0;
  assign _T_4775 = rvx_signal_162[13];
  assign _GEN_3243 = {{13'd0}, rvx_signal_096};
  assign _T_4790 = _GEN_3243 << 13;
  assign _GEN_3244 = {{1'd0}, _T_4754};
  assign _T_4794 = _GEN_3244 | _T_4790;
  assign _T_4802 = _T_4234[14];
  assign _T_4806 = ~ _T_4802;
  assign _T_4808 = _T_4806 == 1'h0;
  assign _T_4815 = rvx_signal_162[14];
  assign _GEN_3245 = {{14'd0}, rvx_signal_167};
  assign _T_4830 = _GEN_3245 << 14;
  assign _GEN_3246 = {{1'd0}, _T_4794};
  assign _T_4834 = _GEN_3246 | _T_4830;
  assign _T_4842 = _T_4234[15];
  assign _T_4846 = ~ _T_4842;
  assign _T_4848 = _T_4846 == 1'h0;
  assign _T_4855 = rvx_signal_162[15];
  assign _GEN_3247 = {{15'd0}, rvx_signal_294};
  assign _T_4870 = _GEN_3247 << 15;
  assign _GEN_3248 = {{1'd0}, _T_4834};
  assign _T_4874 = _GEN_3248 | _T_4870;
  assign _T_4882 = _T_4234[16];
  assign _T_4886 = ~ _T_4882;
  assign _T_4888 = _T_4886 == 1'h0;
  assign _T_4895 = rvx_signal_162[16];
  assign _GEN_3249 = {{16'd0}, rvx_signal_371};
  assign _T_4910 = _GEN_3249 << 16;
  assign _GEN_3250 = {{1'd0}, _T_4874};
  assign _T_4914 = _GEN_3250 | _T_4910;
  assign _T_4922 = _T_4234[17];
  assign _T_4926 = ~ _T_4922;
  assign _T_4928 = _T_4926 == 1'h0;
  assign _T_4935 = rvx_signal_162[17];
  assign _GEN_3251 = {{17'd0}, rvx_signal_103};
  assign _T_4950 = _GEN_3251 << 17;
  assign _GEN_3252 = {{1'd0}, _T_4914};
  assign _T_4954 = _GEN_3252 | _T_4950;
  assign _T_4962 = _T_4234[18];
  assign _T_4966 = ~ _T_4962;
  assign _T_4968 = _T_4966 == 1'h0;
  assign _T_4975 = rvx_signal_162[18];
  assign _GEN_3253 = {{18'd0}, rvx_signal_019};
  assign _T_4990 = _GEN_3253 << 18;
  assign _GEN_3254 = {{1'd0}, _T_4954};
  assign _T_4994 = _GEN_3254 | _T_4990;
  assign _T_5002 = _T_4234[19];
  assign _T_5006 = ~ _T_5002;
  assign _T_5008 = _T_5006 == 1'h0;
  assign _T_5015 = rvx_signal_162[19];
  assign _GEN_3255 = {{19'd0}, rvx_signal_080};
  assign _T_5030 = _GEN_3255 << 19;
  assign _GEN_3256 = {{1'd0}, _T_4994};
  assign _T_5034 = _GEN_3256 | _T_5030;
  assign _T_5042 = _T_4234[20];
  assign _T_5046 = ~ _T_5042;
  assign _T_5048 = _T_5046 == 1'h0;
  assign _T_5055 = rvx_signal_162[20];
  assign _GEN_3257 = {{20'd0}, rvx_signal_239};
  assign _T_5070 = _GEN_3257 << 20;
  assign _GEN_3258 = {{1'd0}, _T_5034};
  assign _T_5074 = _GEN_3258 | _T_5070;
  assign _T_5082 = _T_4234[21];
  assign _T_5086 = ~ _T_5082;
  assign _T_5088 = _T_5086 == 1'h0;
  assign _T_5095 = rvx_signal_162[21];
  assign _GEN_3259 = {{21'd0}, rvx_signal_124};
  assign _T_5110 = _GEN_3259 << 21;
  assign _GEN_3260 = {{1'd0}, _T_5074};
  assign _T_5114 = _GEN_3260 | _T_5110;
  assign _T_5122 = _T_4234[22];
  assign _T_5126 = ~ _T_5122;
  assign _T_5128 = _T_5126 == 1'h0;
  assign _T_5135 = rvx_signal_162[22];
  assign _GEN_3261 = {{22'd0}, rvx_signal_222};
  assign _T_5150 = _GEN_3261 << 22;
  assign _GEN_3262 = {{1'd0}, _T_5114};
  assign _T_5154 = _GEN_3262 | _T_5150;
  assign _T_5162 = _T_4234[23];
  assign _T_5166 = ~ _T_5162;
  assign _T_5168 = _T_5166 == 1'h0;
  assign _T_5175 = rvx_signal_162[23];
  assign _GEN_3263 = {{23'd0}, rvx_signal_306};
  assign _T_5190 = _GEN_3263 << 23;
  assign _GEN_3264 = {{1'd0}, _T_5154};
  assign _T_5194 = _GEN_3264 | _T_5190;
  assign _T_5202 = _T_4234[24];
  assign _T_5206 = ~ _T_5202;
  assign _T_5208 = _T_5206 == 1'h0;
  assign _T_5215 = rvx_signal_162[24];
  assign _GEN_3265 = {{24'd0}, rvx_signal_238};
  assign _T_5230 = _GEN_3265 << 24;
  assign _GEN_3266 = {{1'd0}, _T_5194};
  assign _T_5234 = _GEN_3266 | _T_5230;
  assign _T_5242 = _T_4234[25];
  assign _T_5246 = ~ _T_5242;
  assign _T_5248 = _T_5246 == 1'h0;
  assign _T_5255 = rvx_signal_162[25];
  assign _GEN_3267 = {{25'd0}, rvx_signal_011};
  assign _T_5270 = _GEN_3267 << 25;
  assign _GEN_3268 = {{1'd0}, _T_5234};
  assign _T_5274 = _GEN_3268 | _T_5270;
  assign _T_5282 = _T_4234[26];
  assign _T_5286 = ~ _T_5282;
  assign _T_5288 = _T_5286 == 1'h0;
  assign _T_5295 = rvx_signal_162[26];
  assign _GEN_3269 = {{26'd0}, rvx_signal_029};
  assign _T_5310 = _GEN_3269 << 26;
  assign _GEN_3270 = {{1'd0}, _T_5274};
  assign _T_5314 = _GEN_3270 | _T_5310;
  assign _T_5322 = _T_4234[27];
  assign _T_5326 = ~ _T_5322;
  assign _T_5328 = _T_5326 == 1'h0;
  assign _T_5335 = rvx_signal_162[27];
  assign _GEN_3271 = {{27'd0}, rvx_signal_166};
  assign _T_5350 = _GEN_3271 << 27;
  assign _GEN_3272 = {{1'd0}, _T_5314};
  assign _T_5354 = _GEN_3272 | _T_5350;
  assign _T_5362 = _T_4234[28];
  assign _T_5366 = ~ _T_5362;
  assign _T_5368 = _T_5366 == 1'h0;
  assign _T_5375 = rvx_signal_162[28];
  assign _GEN_3273 = {{28'd0}, rvx_signal_228};
  assign _T_5390 = _GEN_3273 << 28;
  assign _GEN_3274 = {{1'd0}, _T_5354};
  assign _T_5394 = _GEN_3274 | _T_5390;
  assign _T_5402 = _T_4234[29];
  assign _T_5406 = ~ _T_5402;
  assign _T_5408 = _T_5406 == 1'h0;
  assign _T_5415 = rvx_signal_162[29];
  assign _GEN_3275 = {{29'd0}, rvx_signal_183};
  assign _T_5430 = _GEN_3275 << 29;
  assign _GEN_3276 = {{1'd0}, _T_5394};
  assign _T_5434 = _GEN_3276 | _T_5430;
  assign _T_5442 = _T_4234[30];
  assign _T_5446 = ~ _T_5442;
  assign _T_5448 = _T_5446 == 1'h0;
  assign _T_5455 = rvx_signal_162[30];
  assign _GEN_3277 = {{30'd0}, rvx_signal_253};
  assign _T_5470 = _GEN_3277 << 30;
  assign _GEN_3278 = {{1'd0}, _T_5434};
  assign _T_5474 = _GEN_3278 | _T_5470;
  assign _T_5482 = _T_4234[31];
  assign _T_5486 = ~ _T_5482;
  assign _T_5488 = _T_5486 == 1'h0;
  assign _T_5495 = rvx_signal_162[31];
  assign _GEN_3279 = {{31'd0}, rvx_signal_033};
  assign _T_5510 = _GEN_3279 << 31;
  assign _GEN_3280 = {{1'd0}, _T_5474};
  assign _T_5514 = _GEN_3280 | _T_5510;
  assign _T_5524 = _T_4234 != 32'h0;
  assign _T_5526 = ~ _T_4234;
  assign _T_5528 = _T_5526 == 32'h0;
  assign _T_5535 = rvx_signal_162;
  assign _T_5574 = _T_3573_33 & _T_5528;
  assign _GEN_41 = _T_5574 ? _T_5535 : {{29'd0}, rvx_signal_117};
  assign _T_5593 = {{29'd0}, rvx_signal_117};
  assign _T_5614 = _T_3573_34 & _T_5528;
  assign _GEN_42 = _T_5614 ? _T_5535 : {{29'd0}, rvx_signal_395};
  assign _T_5633 = {{29'd0}, rvx_signal_395};
  assign _T_5654 = _T_3573_35 & _T_5528;
  assign _GEN_43 = _T_5654 ? _T_5535 : {{29'd0}, rvx_signal_097};
  assign _T_5673 = {{29'd0}, rvx_signal_097};
  assign _T_5694 = _T_3573_36 & _T_5528;
  assign _GEN_44 = _T_5694 ? _T_5535 : {{29'd0}, rvx_signal_267};
  assign _T_5713 = {{29'd0}, rvx_signal_267};
  assign _T_5734 = _T_3573_37 & _T_5528;
  assign _GEN_45 = _T_5734 ? _T_5535 : {{29'd0}, rvx_signal_025};
  assign _T_5753 = {{29'd0}, rvx_signal_025};
  assign _T_5774 = _T_3573_38 & _T_5528;
  assign _GEN_46 = _T_5774 ? _T_5535 : {{29'd0}, rvx_signal_266};
  assign _T_5793 = {{29'd0}, rvx_signal_266};
  assign _T_5814 = _T_3573_39 & _T_4248;
  assign _GEN_47 = _T_5814 ? _T_4255 : rvx_signal_408;
  assign _T_5854 = _T_3573_40 & _T_5528;
  assign _GEN_48 = _T_5854 ? _T_5535 : {{29'd0}, rvx_signal_359};
  assign _T_5873 = {{29'd0}, rvx_signal_359};
  assign _T_5890 = _T_3466_41 & _T_5524;
  assign _T_5894 = _T_3573_41 & _T_5528;
  assign _T_5897 = _T_5535[5:0];
  assign _T_5898 = rvx_signal_120 == _T_5897;
  assign _T_5900 = _T_5898 | rvx_port_41;
  assign _T_5902 = _T_5900 == 1'h0;
  assign _GEN_49 = 6'h1 == rvx_signal_120 ? rvx_signal_099 : 1'h0;
  assign _GEN_50 = 6'h2 == rvx_signal_120 ? rvx_signal_369 : _GEN_49;
  assign _GEN_51 = 6'h3 == rvx_signal_120 ? rvx_signal_221 : _GEN_50;
  assign _GEN_52 = 6'h4 == rvx_signal_120 ? rvx_signal_224 : _GEN_51;
  assign _GEN_53 = 6'h5 == rvx_signal_120 ? rvx_signal_066 : _GEN_52;
  assign _GEN_54 = 6'h6 == rvx_signal_120 ? rvx_signal_111 : _GEN_53;
  assign _GEN_55 = 6'h7 == rvx_signal_120 ? rvx_signal_179 : _GEN_54;
  assign _GEN_56 = 6'h8 == rvx_signal_120 ? rvx_signal_050 : _GEN_55;
  assign _GEN_57 = 6'h9 == rvx_signal_120 ? rvx_signal_215 : _GEN_56;
  assign _GEN_58 = 6'ha == rvx_signal_120 ? rvx_signal_386 : _GEN_57;
  assign _GEN_59 = 6'hb == rvx_signal_120 ? rvx_signal_450 : _GEN_58;
  assign _GEN_60 = 6'hc == rvx_signal_120 ? rvx_signal_399 : _GEN_59;
  assign _GEN_61 = 6'hd == rvx_signal_120 ? rvx_signal_067 : _GEN_60;
  assign _GEN_62 = 6'he == rvx_signal_120 ? rvx_signal_350 : _GEN_61;
  assign _GEN_63 = 6'hf == rvx_signal_120 ? rvx_signal_265 : _GEN_62;
  assign _GEN_64 = 6'h10 == rvx_signal_120 ? rvx_signal_304 : _GEN_63;
  assign _GEN_65 = 6'h11 == rvx_signal_120 ? rvx_signal_058 : _GEN_64;
  assign _GEN_66 = 6'h12 == rvx_signal_120 ? rvx_signal_433 : _GEN_65;
  assign _GEN_67 = 6'h13 == rvx_signal_120 ? rvx_signal_465 : _GEN_66;
  assign _GEN_68 = 6'h14 == rvx_signal_120 ? rvx_signal_197 : _GEN_67;
  assign _GEN_69 = 6'h15 == rvx_signal_120 ? rvx_signal_358 : _GEN_68;
  assign _GEN_70 = 6'h16 == rvx_signal_120 ? rvx_signal_436 : _GEN_69;
  assign _GEN_71 = 6'h17 == rvx_signal_120 ? rvx_signal_001 : _GEN_70;
  assign _GEN_72 = 6'h18 == rvx_signal_120 ? rvx_signal_131 : _GEN_71;
  assign _GEN_73 = 6'h19 == rvx_signal_120 ? rvx_signal_410 : _GEN_72;
  assign _GEN_74 = 6'h1a == rvx_signal_120 ? rvx_signal_137 : _GEN_73;
  assign _GEN_75 = 6'h1b == rvx_signal_120 ? rvx_signal_178 : _GEN_74;
  assign _GEN_76 = 6'h1c == rvx_signal_120 ? rvx_signal_052 : _GEN_75;
  assign _GEN_77 = 6'h1d == rvx_signal_120 ? rvx_signal_423 : _GEN_76;
  assign _GEN_78 = 6'h1e == rvx_signal_120 ? rvx_signal_462 : _GEN_77;
  assign _GEN_79 = 6'h1f == rvx_signal_120 ? rvx_signal_475 : _GEN_78;
  assign _GEN_80 = 6'h20 == rvx_signal_120 ? rvx_signal_408 : _GEN_79;
  assign _T_5906 = _T_5894 & _GEN_0;
  assign _T_5923 = {{26'd0}, rvx_signal_153};
  assign _T_5944 = _T_3573_42 & _T_5528;
  assign _GEN_81 = _T_5944 ? _T_5535 : {{29'd0}, rvx_signal_243};
  assign _T_5963 = {{29'd0}, rvx_signal_243};
  assign _T_5984 = _T_3573_43 & _T_5528;
  assign _GEN_82 = _T_5984 ? _T_5535 : {{29'd0}, rvx_signal_116};
  assign _T_6003 = {{29'd0}, rvx_signal_116};
  assign _T_6024 = _T_3573_44 & _T_5528;
  assign _GEN_83 = _T_6024 ? _T_5535 : {{29'd0}, rvx_signal_430};
  assign _T_6043 = {{29'd0}, rvx_signal_430};
  assign _T_6064 = _T_3573_45 & _T_5528;
  assign _GEN_84 = _T_6064 ? _T_5535 : {{29'd0}, rvx_signal_444};
  assign _T_6083 = {{29'd0}, rvx_signal_444};
  assign _T_6104 = _T_3573_46 & _T_5528;
  assign _GEN_85 = _T_6104 ? _T_5535 : {{29'd0}, rvx_signal_002};
  assign _T_6123 = {{29'd0}, rvx_signal_002};
  assign _T_6144 = _T_3573_47 & _T_5528;
  assign _GEN_86 = _T_6144 ? _T_5535 : {{29'd0}, rvx_signal_145};
  assign _T_6163 = {{29'd0}, rvx_signal_145};
  assign _T_6184 = _T_3573_48 & _T_5528;
  assign _GEN_87 = _T_6184 ? _T_5535 : {{29'd0}, rvx_signal_057};
  assign _T_6203 = {{29'd0}, rvx_signal_057};
  assign _T_6224 = _T_3573_49 & _T_5528;
  assign _GEN_88 = _T_6224 ? _T_5535 : {{29'd0}, rvx_signal_032};
  assign _T_6243 = {{29'd0}, rvx_signal_032};
  assign _T_6264 = _T_3573_50 & _T_5528;
  assign _GEN_89 = _T_6264 ? _T_5535 : {{29'd0}, rvx_signal_245};
  assign _T_6283 = {{29'd0}, rvx_signal_245};
  assign _T_6304 = _T_3573_51 & _T_5528;
  assign _GEN_90 = _T_6304 ? _T_5535 : {{29'd0}, rvx_signal_435};
  assign _T_6323 = {{29'd0}, rvx_signal_435};
  assign _T_6384 = _T_3573_53 & _T_4288;
  assign _GEN_92 = _T_6384 ? _T_4295 : rvx_signal_099;
  assign _GEN_3281 = {{1'd0}, rvx_signal_099};
  assign _T_6400 = _GEN_3281 << 1;
  assign _T_6424 = _T_3573_54 & _T_4328;
  assign _GEN_93 = _T_6424 ? _T_4335 : rvx_signal_369;
  assign _GEN_3282 = {{2'd0}, rvx_signal_369};
  assign _T_6440 = _GEN_3282 << 2;
  assign _GEN_3283 = {{1'd0}, _T_6400};
  assign _T_6444 = _GEN_3283 | _T_6440;
  assign _T_6464 = _T_3573_55 & _T_4368;
  assign _GEN_94 = _T_6464 ? _T_4375 : rvx_signal_221;
  assign _GEN_3284 = {{3'd0}, rvx_signal_221};
  assign _T_6480 = _GEN_3284 << 3;
  assign _GEN_3285 = {{1'd0}, _T_6444};
  assign _T_6484 = _GEN_3285 | _T_6480;
  assign _T_6504 = _T_3573_56 & _T_4408;
  assign _GEN_95 = _T_6504 ? _T_4415 : rvx_signal_224;
  assign _GEN_3286 = {{4'd0}, rvx_signal_224};
  assign _T_6520 = _GEN_3286 << 4;
  assign _GEN_3287 = {{1'd0}, _T_6484};
  assign _T_6524 = _GEN_3287 | _T_6520;
  assign _T_6544 = _T_3573_57 & _T_4448;
  assign _GEN_96 = _T_6544 ? _T_4455 : rvx_signal_066;
  assign _GEN_3288 = {{5'd0}, rvx_signal_066};
  assign _T_6560 = _GEN_3288 << 5;
  assign _GEN_3289 = {{1'd0}, _T_6524};
  assign _T_6564 = _GEN_3289 | _T_6560;
  assign _T_6584 = _T_3573_58 & _T_4488;
  assign _GEN_97 = _T_6584 ? _T_4495 : rvx_signal_111;
  assign _GEN_3290 = {{6'd0}, rvx_signal_111};
  assign _T_6600 = _GEN_3290 << 6;
  assign _GEN_3291 = {{1'd0}, _T_6564};
  assign _T_6604 = _GEN_3291 | _T_6600;
  assign _T_6624 = _T_3573_59 & _T_4528;
  assign _GEN_98 = _T_6624 ? _T_4535 : rvx_signal_179;
  assign _GEN_3292 = {{7'd0}, rvx_signal_179};
  assign _T_6640 = _GEN_3292 << 7;
  assign _GEN_3293 = {{1'd0}, _T_6604};
  assign _T_6644 = _GEN_3293 | _T_6640;
  assign _T_6664 = _T_3573_60 & _T_4568;
  assign _GEN_99 = _T_6664 ? _T_4575 : rvx_signal_050;
  assign _GEN_3294 = {{8'd0}, rvx_signal_050};
  assign _T_6680 = _GEN_3294 << 8;
  assign _GEN_3295 = {{1'd0}, _T_6644};
  assign _T_6684 = _GEN_3295 | _T_6680;
  assign _T_6704 = _T_3573_61 & _T_4608;
  assign _GEN_100 = _T_6704 ? _T_4615 : rvx_signal_215;
  assign _GEN_3296 = {{9'd0}, rvx_signal_215};
  assign _T_6720 = _GEN_3296 << 9;
  assign _GEN_3297 = {{1'd0}, _T_6684};
  assign _T_6724 = _GEN_3297 | _T_6720;
  assign _T_6744 = _T_3573_62 & _T_4648;
  assign _GEN_101 = _T_6744 ? _T_4655 : rvx_signal_386;
  assign _GEN_3298 = {{10'd0}, rvx_signal_386};
  assign _T_6760 = _GEN_3298 << 10;
  assign _GEN_3299 = {{1'd0}, _T_6724};
  assign _T_6764 = _GEN_3299 | _T_6760;
  assign _T_6784 = _T_3573_63 & _T_4688;
  assign _GEN_102 = _T_6784 ? _T_4695 : rvx_signal_450;
  assign _GEN_3300 = {{11'd0}, rvx_signal_450};
  assign _T_6800 = _GEN_3300 << 11;
  assign _GEN_3301 = {{1'd0}, _T_6764};
  assign _T_6804 = _GEN_3301 | _T_6800;
  assign _T_6824 = _T_3573_64 & _T_4728;
  assign _GEN_103 = _T_6824 ? _T_4735 : rvx_signal_399;
  assign _GEN_3302 = {{12'd0}, rvx_signal_399};
  assign _T_6840 = _GEN_3302 << 12;
  assign _GEN_3303 = {{1'd0}, _T_6804};
  assign _T_6844 = _GEN_3303 | _T_6840;
  assign _T_6864 = _T_3573_65 & _T_4768;
  assign _GEN_104 = _T_6864 ? _T_4775 : rvx_signal_067;
  assign _GEN_3304 = {{13'd0}, rvx_signal_067};
  assign _T_6880 = _GEN_3304 << 13;
  assign _GEN_3305 = {{1'd0}, _T_6844};
  assign _T_6884 = _GEN_3305 | _T_6880;
  assign _T_6904 = _T_3573_66 & _T_4808;
  assign _GEN_105 = _T_6904 ? _T_4815 : rvx_signal_350;
  assign _GEN_3306 = {{14'd0}, rvx_signal_350};
  assign _T_6920 = _GEN_3306 << 14;
  assign _GEN_3307 = {{1'd0}, _T_6884};
  assign _T_6924 = _GEN_3307 | _T_6920;
  assign _T_6944 = _T_3573_67 & _T_4848;
  assign _GEN_106 = _T_6944 ? _T_4855 : rvx_signal_265;
  assign _GEN_3308 = {{15'd0}, rvx_signal_265};
  assign _T_6960 = _GEN_3308 << 15;
  assign _GEN_3309 = {{1'd0}, _T_6924};
  assign _T_6964 = _GEN_3309 | _T_6960;
  assign _T_6984 = _T_3573_68 & _T_4888;
  assign _GEN_107 = _T_6984 ? _T_4895 : rvx_signal_304;
  assign _GEN_3310 = {{16'd0}, rvx_signal_304};
  assign _T_7000 = _GEN_3310 << 16;
  assign _GEN_3311 = {{1'd0}, _T_6964};
  assign _T_7004 = _GEN_3311 | _T_7000;
  assign _T_7024 = _T_3573_69 & _T_4928;
  assign _GEN_108 = _T_7024 ? _T_4935 : rvx_signal_058;
  assign _GEN_3312 = {{17'd0}, rvx_signal_058};
  assign _T_7040 = _GEN_3312 << 17;
  assign _GEN_3313 = {{1'd0}, _T_7004};
  assign _T_7044 = _GEN_3313 | _T_7040;
  assign _T_7064 = _T_3573_70 & _T_4968;
  assign _GEN_109 = _T_7064 ? _T_4975 : rvx_signal_433;
  assign _GEN_3314 = {{18'd0}, rvx_signal_433};
  assign _T_7080 = _GEN_3314 << 18;
  assign _GEN_3315 = {{1'd0}, _T_7044};
  assign _T_7084 = _GEN_3315 | _T_7080;
  assign _T_7104 = _T_3573_71 & _T_5008;
  assign _GEN_110 = _T_7104 ? _T_5015 : rvx_signal_465;
  assign _GEN_3316 = {{19'd0}, rvx_signal_465};
  assign _T_7120 = _GEN_3316 << 19;
  assign _GEN_3317 = {{1'd0}, _T_7084};
  assign _T_7124 = _GEN_3317 | _T_7120;
  assign _T_7144 = _T_3573_72 & _T_5048;
  assign _GEN_111 = _T_7144 ? _T_5055 : rvx_signal_197;
  assign _GEN_3318 = {{20'd0}, rvx_signal_197};
  assign _T_7160 = _GEN_3318 << 20;
  assign _GEN_3319 = {{1'd0}, _T_7124};
  assign _T_7164 = _GEN_3319 | _T_7160;
  assign _T_7184 = _T_3573_73 & _T_5088;
  assign _GEN_112 = _T_7184 ? _T_5095 : rvx_signal_358;
  assign _GEN_3320 = {{21'd0}, rvx_signal_358};
  assign _T_7200 = _GEN_3320 << 21;
  assign _GEN_3321 = {{1'd0}, _T_7164};
  assign _T_7204 = _GEN_3321 | _T_7200;
  assign _T_7224 = _T_3573_74 & _T_5128;
  assign _GEN_113 = _T_7224 ? _T_5135 : rvx_signal_436;
  assign _GEN_3322 = {{22'd0}, rvx_signal_436};
  assign _T_7240 = _GEN_3322 << 22;
  assign _GEN_3323 = {{1'd0}, _T_7204};
  assign _T_7244 = _GEN_3323 | _T_7240;
  assign _T_7264 = _T_3573_75 & _T_5168;
  assign _GEN_114 = _T_7264 ? _T_5175 : rvx_signal_001;
  assign _GEN_3324 = {{23'd0}, rvx_signal_001};
  assign _T_7280 = _GEN_3324 << 23;
  assign _GEN_3325 = {{1'd0}, _T_7244};
  assign _T_7284 = _GEN_3325 | _T_7280;
  assign _T_7304 = _T_3573_76 & _T_5208;
  assign _GEN_115 = _T_7304 ? _T_5215 : rvx_signal_131;
  assign _GEN_3326 = {{24'd0}, rvx_signal_131};
  assign _T_7320 = _GEN_3326 << 24;
  assign _GEN_3327 = {{1'd0}, _T_7284};
  assign _T_7324 = _GEN_3327 | _T_7320;
  assign _T_7344 = _T_3573_77 & _T_5248;
  assign _GEN_116 = _T_7344 ? _T_5255 : rvx_signal_410;
  assign _GEN_3328 = {{25'd0}, rvx_signal_410};
  assign _T_7360 = _GEN_3328 << 25;
  assign _GEN_3329 = {{1'd0}, _T_7324};
  assign _T_7364 = _GEN_3329 | _T_7360;
  assign _T_7384 = _T_3573_78 & _T_5288;
  assign _GEN_117 = _T_7384 ? _T_5295 : rvx_signal_137;
  assign _GEN_3330 = {{26'd0}, rvx_signal_137};
  assign _T_7400 = _GEN_3330 << 26;
  assign _GEN_3331 = {{1'd0}, _T_7364};
  assign _T_7404 = _GEN_3331 | _T_7400;
  assign _T_7424 = _T_3573_79 & _T_5328;
  assign _GEN_118 = _T_7424 ? _T_5335 : rvx_signal_178;
  assign _GEN_3332 = {{27'd0}, rvx_signal_178};
  assign _T_7440 = _GEN_3332 << 27;
  assign _GEN_3333 = {{1'd0}, _T_7404};
  assign _T_7444 = _GEN_3333 | _T_7440;
  assign _T_7464 = _T_3573_80 & _T_5368;
  assign _GEN_119 = _T_7464 ? _T_5375 : rvx_signal_052;
  assign _GEN_3334 = {{28'd0}, rvx_signal_052};
  assign _T_7480 = _GEN_3334 << 28;
  assign _GEN_3335 = {{1'd0}, _T_7444};
  assign _T_7484 = _GEN_3335 | _T_7480;
  assign _T_7504 = _T_3573_81 & _T_5408;
  assign _GEN_120 = _T_7504 ? _T_5415 : rvx_signal_423;
  assign _GEN_3336 = {{29'd0}, rvx_signal_423};
  assign _T_7520 = _GEN_3336 << 29;
  assign _GEN_3337 = {{1'd0}, _T_7484};
  assign _T_7524 = _GEN_3337 | _T_7520;
  assign _T_7544 = _T_3573_82 & _T_5448;
  assign _GEN_121 = _T_7544 ? _T_5455 : rvx_signal_462;
  assign _GEN_3338 = {{30'd0}, rvx_signal_462};
  assign _T_7560 = _GEN_3338 << 30;
  assign _GEN_3339 = {{1'd0}, _T_7524};
  assign _T_7564 = _GEN_3339 | _T_7560;
  assign _T_7584 = _T_3573_83 & _T_5488;
  assign _GEN_122 = _T_7584 ? _T_5495 : rvx_signal_475;
  assign _GEN_3340 = {{31'd0}, rvx_signal_475};
  assign _T_7600 = _GEN_3340 << 31;
  assign _GEN_3341 = {{1'd0}, _T_7564};
  assign _T_7604 = _GEN_3341 | _T_7600;
  assign _T_7624 = _T_3573_84 & _T_5528;
  assign _GEN_123 = _T_7624 ? _T_5535 : {{29'd0}, rvx_signal_088};
  assign _T_7643 = {{29'd0}, rvx_signal_088};
  assign _T_7664 = _T_3573_85 & _T_5528;
  assign _GEN_124 = _T_7664 ? _T_5535 : {{29'd0}, rvx_signal_400};
  assign _T_7683 = {{29'd0}, rvx_signal_400};
  assign _T_7704 = _T_3573_86 & _T_5528;
  assign _GEN_125 = _T_7704 ? _T_5535 : {{29'd0}, rvx_signal_023};
  assign _T_7723 = {{29'd0}, rvx_signal_023};
  assign _T_7744 = _T_3573_87 & _T_5528;
  assign _GEN_126 = _T_7744 ? _T_5535 : {{29'd0}, rvx_signal_415};
  assign _T_7763 = {{29'd0}, rvx_signal_415};
  assign _T_7784 = _T_3573_88 & _T_5528;
  assign _GEN_127 = _T_7784 ? _T_5535 : {{29'd0}, rvx_signal_311};
  assign _T_7803 = {{29'd0}, rvx_signal_311};
  assign _T_7864 = _T_3573_90 & _T_5528;
  assign _GEN_128 = _T_7864 ? _T_5535 : {{29'd0}, rvx_signal_114};
  assign _T_7883 = {{29'd0}, rvx_signal_114};
  assign _T_7904 = _T_3573_91 & _T_5528;
  assign _GEN_129 = _T_7904 ? _T_5535 : {{29'd0}, rvx_signal_008};
  assign _T_7923 = {{29'd0}, rvx_signal_008};
  assign _T_7944 = _T_3573_92 & _T_5528;
  assign _GEN_130 = _T_7944 ? _T_5535 : {{29'd0}, rvx_signal_300};
  assign _T_7963 = {{29'd0}, rvx_signal_300};
  assign _T_7984 = _T_3573_93 & _T_5528;
  assign _GEN_131 = _T_7984 ? _T_5535 : {{29'd0}, rvx_signal_140};
  assign _T_8003 = {{29'd0}, rvx_signal_140};
  assign _T_8024 = _T_3573_94 & _T_5528;
  assign _GEN_132 = _T_8024 ? _T_5535 : {{29'd0}, rvx_signal_248};
  assign _T_8043 = {{29'd0}, rvx_signal_248};
  assign _T_8064 = _T_3573_95 & _T_5528;
  assign _GEN_133 = _T_8064 ? _T_5535 : {{29'd0}, rvx_signal_234};
  assign _T_8083 = {{29'd0}, rvx_signal_234};
  assign _T_8104 = _T_3573_96 & _T_5528;
  assign _GEN_134 = _T_8104 ? _T_5535 : {{29'd0}, rvx_signal_289};
  assign _T_8123 = {{29'd0}, rvx_signal_289};
  assign _T_8144 = _T_3573_97 & _T_5528;
  assign _GEN_135 = _T_8144 ? _T_5535 : {{29'd0}, rvx_signal_332};
  assign _T_8163 = {{29'd0}, rvx_signal_332};
  assign _T_8184 = _T_3573_98 & _T_5528;
  assign _GEN_136 = _T_8184 ? _T_5535 : {{29'd0}, rvx_signal_172};
  assign _T_8203 = {{29'd0}, rvx_signal_172};
  assign _T_8224 = _T_3573_99 & _T_5528;
  assign _GEN_137 = _T_8224 ? _T_5535 : {{29'd0}, rvx_signal_089};
  assign _T_8243 = {{29'd0}, rvx_signal_089};
  assign _T_8264 = _T_3573_100 & _T_5528;
  assign _GEN_138 = _T_8264 ? _T_5535 : {{29'd0}, rvx_signal_418};
  assign _T_8283 = {{29'd0}, rvx_signal_418};
  assign _T_8317 = rvx_signal_060[0];
  assign _T_8318 = rvx_signal_060[1];
  assign _T_8319 = rvx_signal_060[2];
  assign _T_8320 = rvx_signal_060[3];
  assign _T_8321 = rvx_signal_060[4];
  assign _T_8322 = rvx_signal_060[5];
  assign _T_8327 = rvx_signal_060[10];
  assign _T_8328 = rvx_signal_060[11];
  assign _T_8336 = rvx_signal_060[19];
  assign _T_8341 = {_T_8318,_T_8317};
  assign _T_8342 = {_T_8320,_T_8319};
  assign _T_8343 = {_T_8342,_T_8341};
  assign _T_8344 = {_T_8322,_T_8321};
  assign _T_8345 = {_T_8336,_T_8328};
  assign _T_8346 = {_T_8345,_T_8327};
  assign _T_8347 = {_T_8346,_T_8344};
  assign _T_8348 = {_T_8347,_T_8343};
  assign _T_8864 = 512'h1 << _T_8348;
  assign _T_8866 = _T_8864[1];
  assign _T_8867 = _T_8864[2];
  assign _T_8868 = _T_8864[3];
  assign _T_8869 = _T_8864[4];
  assign _T_8870 = _T_8864[5];
  assign _T_8871 = _T_8864[6];
  assign _T_8872 = _T_8864[7];
  assign _T_8873 = _T_8864[8];
  assign _T_8874 = _T_8864[9];
  assign _T_8875 = _T_8864[10];
  assign _T_8876 = _T_8864[11];
  assign _T_8877 = _T_8864[12];
  assign _T_8878 = _T_8864[13];
  assign _T_8879 = _T_8864[14];
  assign _T_8880 = _T_8864[15];
  assign _T_8881 = _T_8864[16];
  assign _T_8882 = _T_8864[17];
  assign _T_8883 = _T_8864[18];
  assign _T_8884 = _T_8864[19];
  assign _T_8885 = _T_8864[20];
  assign _T_8886 = _T_8864[21];
  assign _T_8887 = _T_8864[22];
  assign _T_8888 = _T_8864[23];
  assign _T_8889 = _T_8864[24];
  assign _T_8890 = _T_8864[25];
  assign _T_8891 = _T_8864[26];
  assign _T_8892 = _T_8864[27];
  assign _T_8893 = _T_8864[28];
  assign _T_8894 = _T_8864[29];
  assign _T_8895 = _T_8864[30];
  assign _T_8896 = _T_8864[31];
  assign _T_8897 = _T_8864[32];
  assign _T_8993 = _T_8864[128];
  assign _T_8994 = _T_8864[129];
  assign _T_9121 = _T_8864[256];
  assign _T_9122 = _T_8864[257];
  assign _T_18609 = rvx_signal_309 & _T_1859_ready;
  assign _T_18610 = _T_18609 & rvx_signal_388;
  assign _T_20669 = _T_18610 & _T_9122;
  assign _T_20670 = _T_20669 & _T_2996;
  assign _T_23226 = rvx_signal_388 == 1'h0;
  assign _T_23227 = _T_18609 & _T_23226;
  assign _T_23238 = _T_23227 & _T_8866;
  assign _T_23239 = _T_23238 & _T_3005;
  assign _T_23246 = _T_23227 & _T_8867;
  assign _T_23247 = _T_23246 & _T_3059;
  assign _T_23254 = _T_23227 & _T_8868;
  assign _T_23255 = _T_23254 & _T_3140;
  assign _T_23262 = _T_23227 & _T_8869;
  assign _T_23263 = _T_23262 & _T_3239;
  assign _T_23270 = _T_23227 & _T_8870;
  assign _T_23271 = _T_23270 & _T_2924;
  assign _T_23278 = _T_23227 & _T_8871;
  assign _T_23279 = _T_23278 & _T_3014;
  assign _T_23286 = _T_23227 & _T_8872;
  assign _T_23287 = _T_23286 & _T_3131;
  assign _T_23294 = _T_23227 & _T_8873;
  assign _T_23295 = _T_23294 & _T_3212;
  assign _T_23302 = _T_23227 & _T_8874;
  assign _T_23303 = _T_23302 & _T_3041;
  assign _T_23310 = _T_23227 & _T_8875;
  assign _T_23311 = _T_23310 & _T_2933;
  assign _T_23318 = _T_23227 & _T_8876;
  assign _T_23319 = _T_23318 & _T_3185;
  assign _T_23326 = _T_23227 & _T_8877;
  assign _T_23327 = _T_23326 & _T_3122;
  assign _T_23334 = _T_23227 & _T_8878;
  assign _T_23335 = _T_23334 & _T_3050;
  assign _T_23342 = _T_23227 & _T_8879;
  assign _T_23343 = _T_23342 & _T_2960;
  assign _T_23350 = _T_23227 & _T_8880;
  assign _T_23351 = _T_23350 & _T_3248;
  assign _T_23358 = _T_23227 & _T_8881;
  assign _T_23359 = _T_23358 & _T_3167;
  assign _T_23366 = _T_23227 & _T_8882;
  assign _T_23367 = _T_23366 & _T_3077;
  assign _T_23374 = _T_23227 & _T_8883;
  assign _T_23375 = _T_23374 & _T_3158;
  assign _T_23382 = _T_23227 & _T_8884;
  assign _T_23383 = _T_23382 & _T_3230;
  assign _T_23390 = _T_23227 & _T_8885;
  assign _T_23391 = _T_23390 & _T_2969;
  assign _T_23398 = _T_23227 & _T_8886;
  assign _T_23399 = _T_23398 & _T_3032;
  assign _T_23406 = _T_23227 & _T_8887;
  assign _T_23407 = _T_23406 & _T_3104;
  assign _T_23414 = _T_23227 & _T_8888;
  assign _T_23415 = _T_23414 & _T_3203;
  assign _T_23422 = _T_23227 & _T_8889;
  assign _T_23423 = _T_23422 & _T_2942;
  assign _T_23430 = _T_23227 & _T_8890;
  assign _T_23431 = _T_23430 & _T_2951;
  assign _T_23438 = _T_23227 & _T_8891;
  assign _T_23439 = _T_23438 & _T_3194;
  assign _T_23446 = _T_23227 & _T_8892;
  assign _T_23447 = _T_23446 & _T_3113;
  assign _T_23454 = _T_23227 & _T_8893;
  assign _T_23455 = _T_23454 & _T_3023;
  assign _T_23462 = _T_23227 & _T_8894;
  assign _T_23463 = _T_23462 & _T_2987;
  assign _T_23470 = _T_23227 & _T_8895;
  assign _T_23471 = _T_23470 & _T_3221;
  assign _T_23478 = _T_23227 & _T_8896;
  assign _T_23479 = _T_23478 & _T_3176;
  assign _T_23486 = _T_23227 & _T_8897;
  assign _T_23487 = _T_23486 & _T_3068;
  assign _T_24254 = _T_23227 & _T_8993;
  assign _T_24255 = _T_24254 & _T_3095;
  assign _T_24262 = _T_23227 & _T_8994;
  assign _T_24263 = _T_24262 & _T_2978;
  assign _T_25278 = _T_23227 & _T_9121;
  assign _T_25279 = _T_25278 & _T_3086;
  assign _T_25286 = _T_23227 & _T_9122;
  assign _T_25287 = _T_25286 & _T_2996;
  assign _T_27850 = rvx_signal_309;
  assign _GEN_2183 = 9'h1 == _T_8348 ? _T_27853_1 : _T_27853_0;
  assign _GEN_2184 = 9'h2 == _T_8348 ? _T_27853_2 : _GEN_2183;
  assign _GEN_2185 = 9'h3 == _T_8348 ? _T_27853_3 : _GEN_2184;
  assign _GEN_2186 = 9'h4 == _T_8348 ? _T_27853_4 : _GEN_2185;
  assign _GEN_2187 = 9'h5 == _T_8348 ? _T_27853_5 : _GEN_2186;
  assign _GEN_2188 = 9'h6 == _T_8348 ? _T_27853_6 : _GEN_2187;
  assign _GEN_2189 = 9'h7 == _T_8348 ? _T_27853_7 : _GEN_2188;
  assign _GEN_2190 = 9'h8 == _T_8348 ? _T_27853_8 : _GEN_2189;
  assign _GEN_2191 = 9'h9 == _T_8348 ? _T_27853_9 : _GEN_2190;
  assign _GEN_2192 = 9'ha == _T_8348 ? _T_27853_10 : _GEN_2191;
  assign _GEN_2193 = 9'hb == _T_8348 ? _T_27853_11 : _GEN_2192;
  assign _GEN_2194 = 9'hc == _T_8348 ? _T_27853_12 : _GEN_2193;
  assign _GEN_2195 = 9'hd == _T_8348 ? _T_27853_13 : _GEN_2194;
  assign _GEN_2196 = 9'he == _T_8348 ? _T_27853_14 : _GEN_2195;
  assign _GEN_2197 = 9'hf == _T_8348 ? _T_27853_15 : _GEN_2196;
  assign _GEN_2198 = 9'h10 == _T_8348 ? _T_27853_16 : _GEN_2197;
  assign _GEN_2199 = 9'h11 == _T_8348 ? _T_27853_17 : _GEN_2198;
  assign _GEN_2200 = 9'h12 == _T_8348 ? _T_27853_18 : _GEN_2199;
  assign _GEN_2201 = 9'h13 == _T_8348 ? _T_27853_19 : _GEN_2200;
  assign _GEN_2202 = 9'h14 == _T_8348 ? _T_27853_20 : _GEN_2201;
  assign _GEN_2203 = 9'h15 == _T_8348 ? _T_27853_21 : _GEN_2202;
  assign _GEN_2204 = 9'h16 == _T_8348 ? _T_27853_22 : _GEN_2203;
  assign _GEN_2205 = 9'h17 == _T_8348 ? _T_27853_23 : _GEN_2204;
  assign _GEN_2206 = 9'h18 == _T_8348 ? _T_27853_24 : _GEN_2205;
  assign _GEN_2207 = 9'h19 == _T_8348 ? _T_27853_25 : _GEN_2206;
  assign _GEN_2208 = 9'h1a == _T_8348 ? _T_27853_26 : _GEN_2207;
  assign _GEN_2209 = 9'h1b == _T_8348 ? _T_27853_27 : _GEN_2208;
  assign _GEN_2210 = 9'h1c == _T_8348 ? _T_27853_28 : _GEN_2209;
  assign _GEN_2211 = 9'h1d == _T_8348 ? _T_27853_29 : _GEN_2210;
  assign _GEN_2212 = 9'h1e == _T_8348 ? _T_27853_30 : _GEN_2211;
  assign _GEN_2213 = 9'h1f == _T_8348 ? _T_27853_31 : _GEN_2212;
  assign _GEN_2214 = 9'h20 == _T_8348 ? _T_27853_32 : _GEN_2213;
  assign _GEN_2215 = 9'h21 == _T_8348 ? 1'h1 : _GEN_2214;
  assign _GEN_2216 = 9'h22 == _T_8348 ? 1'h1 : _GEN_2215;
  assign _GEN_2217 = 9'h23 == _T_8348 ? 1'h1 : _GEN_2216;
  assign _GEN_2218 = 9'h24 == _T_8348 ? 1'h1 : _GEN_2217;
  assign _GEN_2219 = 9'h25 == _T_8348 ? 1'h1 : _GEN_2218;
  assign _GEN_2220 = 9'h26 == _T_8348 ? 1'h1 : _GEN_2219;
  assign _GEN_2221 = 9'h27 == _T_8348 ? 1'h1 : _GEN_2220;
  assign _GEN_2222 = 9'h28 == _T_8348 ? 1'h1 : _GEN_2221;
  assign _GEN_2223 = 9'h29 == _T_8348 ? 1'h1 : _GEN_2222;
  assign _GEN_2224 = 9'h2a == _T_8348 ? 1'h1 : _GEN_2223;
  assign _GEN_2225 = 9'h2b == _T_8348 ? 1'h1 : _GEN_2224;
  assign _GEN_2226 = 9'h2c == _T_8348 ? 1'h1 : _GEN_2225;
  assign _GEN_2227 = 9'h2d == _T_8348 ? 1'h1 : _GEN_2226;
  assign _GEN_2228 = 9'h2e == _T_8348 ? 1'h1 : _GEN_2227;
  assign _GEN_2229 = 9'h2f == _T_8348 ? 1'h1 : _GEN_2228;
  assign _GEN_2230 = 9'h30 == _T_8348 ? 1'h1 : _GEN_2229;
  assign _GEN_2231 = 9'h31 == _T_8348 ? 1'h1 : _GEN_2230;
  assign _GEN_2232 = 9'h32 == _T_8348 ? 1'h1 : _GEN_2231;
  assign _GEN_2233 = 9'h33 == _T_8348 ? 1'h1 : _GEN_2232;
  assign _GEN_2234 = 9'h34 == _T_8348 ? 1'h1 : _GEN_2233;
  assign _GEN_2235 = 9'h35 == _T_8348 ? 1'h1 : _GEN_2234;
  assign _GEN_2236 = 9'h36 == _T_8348 ? 1'h1 : _GEN_2235;
  assign _GEN_2237 = 9'h37 == _T_8348 ? 1'h1 : _GEN_2236;
  assign _GEN_2238 = 9'h38 == _T_8348 ? 1'h1 : _GEN_2237;
  assign _GEN_2239 = 9'h39 == _T_8348 ? 1'h1 : _GEN_2238;
  assign _GEN_2240 = 9'h3a == _T_8348 ? 1'h1 : _GEN_2239;
  assign _GEN_2241 = 9'h3b == _T_8348 ? 1'h1 : _GEN_2240;
  assign _GEN_2242 = 9'h3c == _T_8348 ? 1'h1 : _GEN_2241;
  assign _GEN_2243 = 9'h3d == _T_8348 ? 1'h1 : _GEN_2242;
  assign _GEN_2244 = 9'h3e == _T_8348 ? 1'h1 : _GEN_2243;
  assign _GEN_2245 = 9'h3f == _T_8348 ? 1'h1 : _GEN_2244;
  assign _GEN_2246 = 9'h40 == _T_8348 ? _T_27853_64 : _GEN_2245;
  assign _GEN_2247 = 9'h41 == _T_8348 ? _T_27853_65 : _GEN_2246;
  assign _GEN_2248 = 9'h42 == _T_8348 ? 1'h1 : _GEN_2247;
  assign _GEN_2249 = 9'h43 == _T_8348 ? 1'h1 : _GEN_2248;
  assign _GEN_2250 = 9'h44 == _T_8348 ? 1'h1 : _GEN_2249;
  assign _GEN_2251 = 9'h45 == _T_8348 ? 1'h1 : _GEN_2250;
  assign _GEN_2252 = 9'h46 == _T_8348 ? 1'h1 : _GEN_2251;
  assign _GEN_2253 = 9'h47 == _T_8348 ? 1'h1 : _GEN_2252;
  assign _GEN_2254 = 9'h48 == _T_8348 ? 1'h1 : _GEN_2253;
  assign _GEN_2255 = 9'h49 == _T_8348 ? 1'h1 : _GEN_2254;
  assign _GEN_2256 = 9'h4a == _T_8348 ? 1'h1 : _GEN_2255;
  assign _GEN_2257 = 9'h4b == _T_8348 ? 1'h1 : _GEN_2256;
  assign _GEN_2258 = 9'h4c == _T_8348 ? 1'h1 : _GEN_2257;
  assign _GEN_2259 = 9'h4d == _T_8348 ? 1'h1 : _GEN_2258;
  assign _GEN_2260 = 9'h4e == _T_8348 ? 1'h1 : _GEN_2259;
  assign _GEN_2261 = 9'h4f == _T_8348 ? 1'h1 : _GEN_2260;
  assign _GEN_2262 = 9'h50 == _T_8348 ? 1'h1 : _GEN_2261;
  assign _GEN_2263 = 9'h51 == _T_8348 ? 1'h1 : _GEN_2262;
  assign _GEN_2264 = 9'h52 == _T_8348 ? 1'h1 : _GEN_2263;
  assign _GEN_2265 = 9'h53 == _T_8348 ? 1'h1 : _GEN_2264;
  assign _GEN_2266 = 9'h54 == _T_8348 ? 1'h1 : _GEN_2265;
  assign _GEN_2267 = 9'h55 == _T_8348 ? 1'h1 : _GEN_2266;
  assign _GEN_2268 = 9'h56 == _T_8348 ? 1'h1 : _GEN_2267;
  assign _GEN_2269 = 9'h57 == _T_8348 ? 1'h1 : _GEN_2268;
  assign _GEN_2270 = 9'h58 == _T_8348 ? 1'h1 : _GEN_2269;
  assign _GEN_2271 = 9'h59 == _T_8348 ? 1'h1 : _GEN_2270;
  assign _GEN_2272 = 9'h5a == _T_8348 ? 1'h1 : _GEN_2271;
  assign _GEN_2273 = 9'h5b == _T_8348 ? 1'h1 : _GEN_2272;
  assign _GEN_2274 = 9'h5c == _T_8348 ? 1'h1 : _GEN_2273;
  assign _GEN_2275 = 9'h5d == _T_8348 ? 1'h1 : _GEN_2274;
  assign _GEN_2276 = 9'h5e == _T_8348 ? 1'h1 : _GEN_2275;
  assign _GEN_2277 = 9'h5f == _T_8348 ? 1'h1 : _GEN_2276;
  assign _GEN_2278 = 9'h60 == _T_8348 ? 1'h1 : _GEN_2277;
  assign _GEN_2279 = 9'h61 == _T_8348 ? 1'h1 : _GEN_2278;
  assign _GEN_2280 = 9'h62 == _T_8348 ? 1'h1 : _GEN_2279;
  assign _GEN_2281 = 9'h63 == _T_8348 ? 1'h1 : _GEN_2280;
  assign _GEN_2282 = 9'h64 == _T_8348 ? 1'h1 : _GEN_2281;
  assign _GEN_2283 = 9'h65 == _T_8348 ? 1'h1 : _GEN_2282;
  assign _GEN_2284 = 9'h66 == _T_8348 ? 1'h1 : _GEN_2283;
  assign _GEN_2285 = 9'h67 == _T_8348 ? 1'h1 : _GEN_2284;
  assign _GEN_2286 = 9'h68 == _T_8348 ? 1'h1 : _GEN_2285;
  assign _GEN_2287 = 9'h69 == _T_8348 ? 1'h1 : _GEN_2286;
  assign _GEN_2288 = 9'h6a == _T_8348 ? 1'h1 : _GEN_2287;
  assign _GEN_2289 = 9'h6b == _T_8348 ? 1'h1 : _GEN_2288;
  assign _GEN_2290 = 9'h6c == _T_8348 ? 1'h1 : _GEN_2289;
  assign _GEN_2291 = 9'h6d == _T_8348 ? 1'h1 : _GEN_2290;
  assign _GEN_2292 = 9'h6e == _T_8348 ? 1'h1 : _GEN_2291;
  assign _GEN_2293 = 9'h6f == _T_8348 ? 1'h1 : _GEN_2292;
  assign _GEN_2294 = 9'h70 == _T_8348 ? 1'h1 : _GEN_2293;
  assign _GEN_2295 = 9'h71 == _T_8348 ? 1'h1 : _GEN_2294;
  assign _GEN_2296 = 9'h72 == _T_8348 ? 1'h1 : _GEN_2295;
  assign _GEN_2297 = 9'h73 == _T_8348 ? 1'h1 : _GEN_2296;
  assign _GEN_2298 = 9'h74 == _T_8348 ? 1'h1 : _GEN_2297;
  assign _GEN_2299 = 9'h75 == _T_8348 ? 1'h1 : _GEN_2298;
  assign _GEN_2300 = 9'h76 == _T_8348 ? 1'h1 : _GEN_2299;
  assign _GEN_2301 = 9'h77 == _T_8348 ? 1'h1 : _GEN_2300;
  assign _GEN_2302 = 9'h78 == _T_8348 ? 1'h1 : _GEN_2301;
  assign _GEN_2303 = 9'h79 == _T_8348 ? 1'h1 : _GEN_2302;
  assign _GEN_2304 = 9'h7a == _T_8348 ? 1'h1 : _GEN_2303;
  assign _GEN_2305 = 9'h7b == _T_8348 ? 1'h1 : _GEN_2304;
  assign _GEN_2306 = 9'h7c == _T_8348 ? 1'h1 : _GEN_2305;
  assign _GEN_2307 = 9'h7d == _T_8348 ? 1'h1 : _GEN_2306;
  assign _GEN_2308 = 9'h7e == _T_8348 ? 1'h1 : _GEN_2307;
  assign _GEN_2309 = 9'h7f == _T_8348 ? 1'h1 : _GEN_2308;
  assign _GEN_2310 = 9'h80 == _T_8348 ? _T_27853_128 : _GEN_2309;
  assign _GEN_2311 = 9'h81 == _T_8348 ? _T_27853_129 : _GEN_2310;
  assign _GEN_2312 = 9'h82 == _T_8348 ? 1'h1 : _GEN_2311;
  assign _GEN_2313 = 9'h83 == _T_8348 ? 1'h1 : _GEN_2312;
  assign _GEN_2314 = 9'h84 == _T_8348 ? 1'h1 : _GEN_2313;
  assign _GEN_2315 = 9'h85 == _T_8348 ? 1'h1 : _GEN_2314;
  assign _GEN_2316 = 9'h86 == _T_8348 ? 1'h1 : _GEN_2315;
  assign _GEN_2317 = 9'h87 == _T_8348 ? 1'h1 : _GEN_2316;
  assign _GEN_2318 = 9'h88 == _T_8348 ? 1'h1 : _GEN_2317;
  assign _GEN_2319 = 9'h89 == _T_8348 ? 1'h1 : _GEN_2318;
  assign _GEN_2320 = 9'h8a == _T_8348 ? 1'h1 : _GEN_2319;
  assign _GEN_2321 = 9'h8b == _T_8348 ? 1'h1 : _GEN_2320;
  assign _GEN_2322 = 9'h8c == _T_8348 ? 1'h1 : _GEN_2321;
  assign _GEN_2323 = 9'h8d == _T_8348 ? 1'h1 : _GEN_2322;
  assign _GEN_2324 = 9'h8e == _T_8348 ? 1'h1 : _GEN_2323;
  assign _GEN_2325 = 9'h8f == _T_8348 ? 1'h1 : _GEN_2324;
  assign _GEN_2326 = 9'h90 == _T_8348 ? 1'h1 : _GEN_2325;
  assign _GEN_2327 = 9'h91 == _T_8348 ? 1'h1 : _GEN_2326;
  assign _GEN_2328 = 9'h92 == _T_8348 ? 1'h1 : _GEN_2327;
  assign _GEN_2329 = 9'h93 == _T_8348 ? 1'h1 : _GEN_2328;
  assign _GEN_2330 = 9'h94 == _T_8348 ? 1'h1 : _GEN_2329;
  assign _GEN_2331 = 9'h95 == _T_8348 ? 1'h1 : _GEN_2330;
  assign _GEN_2332 = 9'h96 == _T_8348 ? 1'h1 : _GEN_2331;
  assign _GEN_2333 = 9'h97 == _T_8348 ? 1'h1 : _GEN_2332;
  assign _GEN_2334 = 9'h98 == _T_8348 ? 1'h1 : _GEN_2333;
  assign _GEN_2335 = 9'h99 == _T_8348 ? 1'h1 : _GEN_2334;
  assign _GEN_2336 = 9'h9a == _T_8348 ? 1'h1 : _GEN_2335;
  assign _GEN_2337 = 9'h9b == _T_8348 ? 1'h1 : _GEN_2336;
  assign _GEN_2338 = 9'h9c == _T_8348 ? 1'h1 : _GEN_2337;
  assign _GEN_2339 = 9'h9d == _T_8348 ? 1'h1 : _GEN_2338;
  assign _GEN_2340 = 9'h9e == _T_8348 ? 1'h1 : _GEN_2339;
  assign _GEN_2341 = 9'h9f == _T_8348 ? 1'h1 : _GEN_2340;
  assign _GEN_2342 = 9'ha0 == _T_8348 ? 1'h1 : _GEN_2341;
  assign _GEN_2343 = 9'ha1 == _T_8348 ? 1'h1 : _GEN_2342;
  assign _GEN_2344 = 9'ha2 == _T_8348 ? 1'h1 : _GEN_2343;
  assign _GEN_2345 = 9'ha3 == _T_8348 ? 1'h1 : _GEN_2344;
  assign _GEN_2346 = 9'ha4 == _T_8348 ? 1'h1 : _GEN_2345;
  assign _GEN_2347 = 9'ha5 == _T_8348 ? 1'h1 : _GEN_2346;
  assign _GEN_2348 = 9'ha6 == _T_8348 ? 1'h1 : _GEN_2347;
  assign _GEN_2349 = 9'ha7 == _T_8348 ? 1'h1 : _GEN_2348;
  assign _GEN_2350 = 9'ha8 == _T_8348 ? 1'h1 : _GEN_2349;
  assign _GEN_2351 = 9'ha9 == _T_8348 ? 1'h1 : _GEN_2350;
  assign _GEN_2352 = 9'haa == _T_8348 ? 1'h1 : _GEN_2351;
  assign _GEN_2353 = 9'hab == _T_8348 ? 1'h1 : _GEN_2352;
  assign _GEN_2354 = 9'hac == _T_8348 ? 1'h1 : _GEN_2353;
  assign _GEN_2355 = 9'had == _T_8348 ? 1'h1 : _GEN_2354;
  assign _GEN_2356 = 9'hae == _T_8348 ? 1'h1 : _GEN_2355;
  assign _GEN_2357 = 9'haf == _T_8348 ? 1'h1 : _GEN_2356;
  assign _GEN_2358 = 9'hb0 == _T_8348 ? 1'h1 : _GEN_2357;
  assign _GEN_2359 = 9'hb1 == _T_8348 ? 1'h1 : _GEN_2358;
  assign _GEN_2360 = 9'hb2 == _T_8348 ? 1'h1 : _GEN_2359;
  assign _GEN_2361 = 9'hb3 == _T_8348 ? 1'h1 : _GEN_2360;
  assign _GEN_2362 = 9'hb4 == _T_8348 ? 1'h1 : _GEN_2361;
  assign _GEN_2363 = 9'hb5 == _T_8348 ? 1'h1 : _GEN_2362;
  assign _GEN_2364 = 9'hb6 == _T_8348 ? 1'h1 : _GEN_2363;
  assign _GEN_2365 = 9'hb7 == _T_8348 ? 1'h1 : _GEN_2364;
  assign _GEN_2366 = 9'hb8 == _T_8348 ? 1'h1 : _GEN_2365;
  assign _GEN_2367 = 9'hb9 == _T_8348 ? 1'h1 : _GEN_2366;
  assign _GEN_2368 = 9'hba == _T_8348 ? 1'h1 : _GEN_2367;
  assign _GEN_2369 = 9'hbb == _T_8348 ? 1'h1 : _GEN_2368;
  assign _GEN_2370 = 9'hbc == _T_8348 ? 1'h1 : _GEN_2369;
  assign _GEN_2371 = 9'hbd == _T_8348 ? 1'h1 : _GEN_2370;
  assign _GEN_2372 = 9'hbe == _T_8348 ? 1'h1 : _GEN_2371;
  assign _GEN_2373 = 9'hbf == _T_8348 ? 1'h1 : _GEN_2372;
  assign _GEN_2374 = 9'hc0 == _T_8348 ? 1'h1 : _GEN_2373;
  assign _GEN_2375 = 9'hc1 == _T_8348 ? 1'h1 : _GEN_2374;
  assign _GEN_2376 = 9'hc2 == _T_8348 ? 1'h1 : _GEN_2375;
  assign _GEN_2377 = 9'hc3 == _T_8348 ? 1'h1 : _GEN_2376;
  assign _GEN_2378 = 9'hc4 == _T_8348 ? 1'h1 : _GEN_2377;
  assign _GEN_2379 = 9'hc5 == _T_8348 ? 1'h1 : _GEN_2378;
  assign _GEN_2380 = 9'hc6 == _T_8348 ? 1'h1 : _GEN_2379;
  assign _GEN_2381 = 9'hc7 == _T_8348 ? 1'h1 : _GEN_2380;
  assign _GEN_2382 = 9'hc8 == _T_8348 ? 1'h1 : _GEN_2381;
  assign _GEN_2383 = 9'hc9 == _T_8348 ? 1'h1 : _GEN_2382;
  assign _GEN_2384 = 9'hca == _T_8348 ? 1'h1 : _GEN_2383;
  assign _GEN_2385 = 9'hcb == _T_8348 ? 1'h1 : _GEN_2384;
  assign _GEN_2386 = 9'hcc == _T_8348 ? 1'h1 : _GEN_2385;
  assign _GEN_2387 = 9'hcd == _T_8348 ? 1'h1 : _GEN_2386;
  assign _GEN_2388 = 9'hce == _T_8348 ? 1'h1 : _GEN_2387;
  assign _GEN_2389 = 9'hcf == _T_8348 ? 1'h1 : _GEN_2388;
  assign _GEN_2390 = 9'hd0 == _T_8348 ? 1'h1 : _GEN_2389;
  assign _GEN_2391 = 9'hd1 == _T_8348 ? 1'h1 : _GEN_2390;
  assign _GEN_2392 = 9'hd2 == _T_8348 ? 1'h1 : _GEN_2391;
  assign _GEN_2393 = 9'hd3 == _T_8348 ? 1'h1 : _GEN_2392;
  assign _GEN_2394 = 9'hd4 == _T_8348 ? 1'h1 : _GEN_2393;
  assign _GEN_2395 = 9'hd5 == _T_8348 ? 1'h1 : _GEN_2394;
  assign _GEN_2396 = 9'hd6 == _T_8348 ? 1'h1 : _GEN_2395;
  assign _GEN_2397 = 9'hd7 == _T_8348 ? 1'h1 : _GEN_2396;
  assign _GEN_2398 = 9'hd8 == _T_8348 ? 1'h1 : _GEN_2397;
  assign _GEN_2399 = 9'hd9 == _T_8348 ? 1'h1 : _GEN_2398;
  assign _GEN_2400 = 9'hda == _T_8348 ? 1'h1 : _GEN_2399;
  assign _GEN_2401 = 9'hdb == _T_8348 ? 1'h1 : _GEN_2400;
  assign _GEN_2402 = 9'hdc == _T_8348 ? 1'h1 : _GEN_2401;
  assign _GEN_2403 = 9'hdd == _T_8348 ? 1'h1 : _GEN_2402;
  assign _GEN_2404 = 9'hde == _T_8348 ? 1'h1 : _GEN_2403;
  assign _GEN_2405 = 9'hdf == _T_8348 ? 1'h1 : _GEN_2404;
  assign _GEN_2406 = 9'he0 == _T_8348 ? 1'h1 : _GEN_2405;
  assign _GEN_2407 = 9'he1 == _T_8348 ? 1'h1 : _GEN_2406;
  assign _GEN_2408 = 9'he2 == _T_8348 ? 1'h1 : _GEN_2407;
  assign _GEN_2409 = 9'he3 == _T_8348 ? 1'h1 : _GEN_2408;
  assign _GEN_2410 = 9'he4 == _T_8348 ? 1'h1 : _GEN_2409;
  assign _GEN_2411 = 9'he5 == _T_8348 ? 1'h1 : _GEN_2410;
  assign _GEN_2412 = 9'he6 == _T_8348 ? 1'h1 : _GEN_2411;
  assign _GEN_2413 = 9'he7 == _T_8348 ? 1'h1 : _GEN_2412;
  assign _GEN_2414 = 9'he8 == _T_8348 ? 1'h1 : _GEN_2413;
  assign _GEN_2415 = 9'he9 == _T_8348 ? 1'h1 : _GEN_2414;
  assign _GEN_2416 = 9'hea == _T_8348 ? 1'h1 : _GEN_2415;
  assign _GEN_2417 = 9'heb == _T_8348 ? 1'h1 : _GEN_2416;
  assign _GEN_2418 = 9'hec == _T_8348 ? 1'h1 : _GEN_2417;
  assign _GEN_2419 = 9'hed == _T_8348 ? 1'h1 : _GEN_2418;
  assign _GEN_2420 = 9'hee == _T_8348 ? 1'h1 : _GEN_2419;
  assign _GEN_2421 = 9'hef == _T_8348 ? 1'h1 : _GEN_2420;
  assign _GEN_2422 = 9'hf0 == _T_8348 ? 1'h1 : _GEN_2421;
  assign _GEN_2423 = 9'hf1 == _T_8348 ? 1'h1 : _GEN_2422;
  assign _GEN_2424 = 9'hf2 == _T_8348 ? 1'h1 : _GEN_2423;
  assign _GEN_2425 = 9'hf3 == _T_8348 ? 1'h1 : _GEN_2424;
  assign _GEN_2426 = 9'hf4 == _T_8348 ? 1'h1 : _GEN_2425;
  assign _GEN_2427 = 9'hf5 == _T_8348 ? 1'h1 : _GEN_2426;
  assign _GEN_2428 = 9'hf6 == _T_8348 ? 1'h1 : _GEN_2427;
  assign _GEN_2429 = 9'hf7 == _T_8348 ? 1'h1 : _GEN_2428;
  assign _GEN_2430 = 9'hf8 == _T_8348 ? 1'h1 : _GEN_2429;
  assign _GEN_2431 = 9'hf9 == _T_8348 ? 1'h1 : _GEN_2430;
  assign _GEN_2432 = 9'hfa == _T_8348 ? 1'h1 : _GEN_2431;
  assign _GEN_2433 = 9'hfb == _T_8348 ? 1'h1 : _GEN_2432;
  assign _GEN_2434 = 9'hfc == _T_8348 ? 1'h1 : _GEN_2433;
  assign _GEN_2435 = 9'hfd == _T_8348 ? 1'h1 : _GEN_2434;
  assign _GEN_2436 = 9'hfe == _T_8348 ? 1'h1 : _GEN_2435;
  assign _GEN_2437 = 9'hff == _T_8348 ? 1'h1 : _GEN_2436;
  assign _GEN_2438 = 9'h100 == _T_8348 ? _T_27853_256 : _GEN_2437;
  assign _GEN_2439 = 9'h101 == _T_8348 ? _T_27853_257 : _GEN_2438;
  assign _GEN_2440 = 9'h102 == _T_8348 ? 1'h1 : _GEN_2439;
  assign _GEN_2441 = 9'h103 == _T_8348 ? 1'h1 : _GEN_2440;
  assign _GEN_2442 = 9'h104 == _T_8348 ? 1'h1 : _GEN_2441;
  assign _GEN_2443 = 9'h105 == _T_8348 ? 1'h1 : _GEN_2442;
  assign _GEN_2444 = 9'h106 == _T_8348 ? 1'h1 : _GEN_2443;
  assign _GEN_2445 = 9'h107 == _T_8348 ? 1'h1 : _GEN_2444;
  assign _GEN_2446 = 9'h108 == _T_8348 ? 1'h1 : _GEN_2445;
  assign _GEN_2447 = 9'h109 == _T_8348 ? 1'h1 : _GEN_2446;
  assign _GEN_2448 = 9'h10a == _T_8348 ? 1'h1 : _GEN_2447;
  assign _GEN_2449 = 9'h10b == _T_8348 ? 1'h1 : _GEN_2448;
  assign _GEN_2450 = 9'h10c == _T_8348 ? 1'h1 : _GEN_2449;
  assign _GEN_2451 = 9'h10d == _T_8348 ? 1'h1 : _GEN_2450;
  assign _GEN_2452 = 9'h10e == _T_8348 ? 1'h1 : _GEN_2451;
  assign _GEN_2453 = 9'h10f == _T_8348 ? 1'h1 : _GEN_2452;
  assign _GEN_2454 = 9'h110 == _T_8348 ? 1'h1 : _GEN_2453;
  assign _GEN_2455 = 9'h111 == _T_8348 ? 1'h1 : _GEN_2454;
  assign _GEN_2456 = 9'h112 == _T_8348 ? 1'h1 : _GEN_2455;
  assign _GEN_2457 = 9'h113 == _T_8348 ? 1'h1 : _GEN_2456;
  assign _GEN_2458 = 9'h114 == _T_8348 ? 1'h1 : _GEN_2457;
  assign _GEN_2459 = 9'h115 == _T_8348 ? 1'h1 : _GEN_2458;
  assign _GEN_2460 = 9'h116 == _T_8348 ? 1'h1 : _GEN_2459;
  assign _GEN_2461 = 9'h117 == _T_8348 ? 1'h1 : _GEN_2460;
  assign _GEN_2462 = 9'h118 == _T_8348 ? 1'h1 : _GEN_2461;
  assign _GEN_2463 = 9'h119 == _T_8348 ? 1'h1 : _GEN_2462;
  assign _GEN_2464 = 9'h11a == _T_8348 ? 1'h1 : _GEN_2463;
  assign _GEN_2465 = 9'h11b == _T_8348 ? 1'h1 : _GEN_2464;
  assign _GEN_2466 = 9'h11c == _T_8348 ? 1'h1 : _GEN_2465;
  assign _GEN_2467 = 9'h11d == _T_8348 ? 1'h1 : _GEN_2466;
  assign _GEN_2468 = 9'h11e == _T_8348 ? 1'h1 : _GEN_2467;
  assign _GEN_2469 = 9'h11f == _T_8348 ? 1'h1 : _GEN_2468;
  assign _GEN_2470 = 9'h120 == _T_8348 ? 1'h1 : _GEN_2469;
  assign _GEN_2471 = 9'h121 == _T_8348 ? 1'h1 : _GEN_2470;
  assign _GEN_2472 = 9'h122 == _T_8348 ? 1'h1 : _GEN_2471;
  assign _GEN_2473 = 9'h123 == _T_8348 ? 1'h1 : _GEN_2472;
  assign _GEN_2474 = 9'h124 == _T_8348 ? 1'h1 : _GEN_2473;
  assign _GEN_2475 = 9'h125 == _T_8348 ? 1'h1 : _GEN_2474;
  assign _GEN_2476 = 9'h126 == _T_8348 ? 1'h1 : _GEN_2475;
  assign _GEN_2477 = 9'h127 == _T_8348 ? 1'h1 : _GEN_2476;
  assign _GEN_2478 = 9'h128 == _T_8348 ? 1'h1 : _GEN_2477;
  assign _GEN_2479 = 9'h129 == _T_8348 ? 1'h1 : _GEN_2478;
  assign _GEN_2480 = 9'h12a == _T_8348 ? 1'h1 : _GEN_2479;
  assign _GEN_2481 = 9'h12b == _T_8348 ? 1'h1 : _GEN_2480;
  assign _GEN_2482 = 9'h12c == _T_8348 ? 1'h1 : _GEN_2481;
  assign _GEN_2483 = 9'h12d == _T_8348 ? 1'h1 : _GEN_2482;
  assign _GEN_2484 = 9'h12e == _T_8348 ? 1'h1 : _GEN_2483;
  assign _GEN_2485 = 9'h12f == _T_8348 ? 1'h1 : _GEN_2484;
  assign _GEN_2486 = 9'h130 == _T_8348 ? 1'h1 : _GEN_2485;
  assign _GEN_2487 = 9'h131 == _T_8348 ? 1'h1 : _GEN_2486;
  assign _GEN_2488 = 9'h132 == _T_8348 ? 1'h1 : _GEN_2487;
  assign _GEN_2489 = 9'h133 == _T_8348 ? 1'h1 : _GEN_2488;
  assign _GEN_2490 = 9'h134 == _T_8348 ? 1'h1 : _GEN_2489;
  assign _GEN_2491 = 9'h135 == _T_8348 ? 1'h1 : _GEN_2490;
  assign _GEN_2492 = 9'h136 == _T_8348 ? 1'h1 : _GEN_2491;
  assign _GEN_2493 = 9'h137 == _T_8348 ? 1'h1 : _GEN_2492;
  assign _GEN_2494 = 9'h138 == _T_8348 ? 1'h1 : _GEN_2493;
  assign _GEN_2495 = 9'h139 == _T_8348 ? 1'h1 : _GEN_2494;
  assign _GEN_2496 = 9'h13a == _T_8348 ? 1'h1 : _GEN_2495;
  assign _GEN_2497 = 9'h13b == _T_8348 ? 1'h1 : _GEN_2496;
  assign _GEN_2498 = 9'h13c == _T_8348 ? 1'h1 : _GEN_2497;
  assign _GEN_2499 = 9'h13d == _T_8348 ? 1'h1 : _GEN_2498;
  assign _GEN_2500 = 9'h13e == _T_8348 ? 1'h1 : _GEN_2499;
  assign _GEN_2501 = 9'h13f == _T_8348 ? 1'h1 : _GEN_2500;
  assign _GEN_2502 = 9'h140 == _T_8348 ? 1'h1 : _GEN_2501;
  assign _GEN_2503 = 9'h141 == _T_8348 ? 1'h1 : _GEN_2502;
  assign _GEN_2504 = 9'h142 == _T_8348 ? 1'h1 : _GEN_2503;
  assign _GEN_2505 = 9'h143 == _T_8348 ? 1'h1 : _GEN_2504;
  assign _GEN_2506 = 9'h144 == _T_8348 ? 1'h1 : _GEN_2505;
  assign _GEN_2507 = 9'h145 == _T_8348 ? 1'h1 : _GEN_2506;
  assign _GEN_2508 = 9'h146 == _T_8348 ? 1'h1 : _GEN_2507;
  assign _GEN_2509 = 9'h147 == _T_8348 ? 1'h1 : _GEN_2508;
  assign _GEN_2510 = 9'h148 == _T_8348 ? 1'h1 : _GEN_2509;
  assign _GEN_2511 = 9'h149 == _T_8348 ? 1'h1 : _GEN_2510;
  assign _GEN_2512 = 9'h14a == _T_8348 ? 1'h1 : _GEN_2511;
  assign _GEN_2513 = 9'h14b == _T_8348 ? 1'h1 : _GEN_2512;
  assign _GEN_2514 = 9'h14c == _T_8348 ? 1'h1 : _GEN_2513;
  assign _GEN_2515 = 9'h14d == _T_8348 ? 1'h1 : _GEN_2514;
  assign _GEN_2516 = 9'h14e == _T_8348 ? 1'h1 : _GEN_2515;
  assign _GEN_2517 = 9'h14f == _T_8348 ? 1'h1 : _GEN_2516;
  assign _GEN_2518 = 9'h150 == _T_8348 ? 1'h1 : _GEN_2517;
  assign _GEN_2519 = 9'h151 == _T_8348 ? 1'h1 : _GEN_2518;
  assign _GEN_2520 = 9'h152 == _T_8348 ? 1'h1 : _GEN_2519;
  assign _GEN_2521 = 9'h153 == _T_8348 ? 1'h1 : _GEN_2520;
  assign _GEN_2522 = 9'h154 == _T_8348 ? 1'h1 : _GEN_2521;
  assign _GEN_2523 = 9'h155 == _T_8348 ? 1'h1 : _GEN_2522;
  assign _GEN_2524 = 9'h156 == _T_8348 ? 1'h1 : _GEN_2523;
  assign _GEN_2525 = 9'h157 == _T_8348 ? 1'h1 : _GEN_2524;
  assign _GEN_2526 = 9'h158 == _T_8348 ? 1'h1 : _GEN_2525;
  assign _GEN_2527 = 9'h159 == _T_8348 ? 1'h1 : _GEN_2526;
  assign _GEN_2528 = 9'h15a == _T_8348 ? 1'h1 : _GEN_2527;
  assign _GEN_2529 = 9'h15b == _T_8348 ? 1'h1 : _GEN_2528;
  assign _GEN_2530 = 9'h15c == _T_8348 ? 1'h1 : _GEN_2529;
  assign _GEN_2531 = 9'h15d == _T_8348 ? 1'h1 : _GEN_2530;
  assign _GEN_2532 = 9'h15e == _T_8348 ? 1'h1 : _GEN_2531;
  assign _GEN_2533 = 9'h15f == _T_8348 ? 1'h1 : _GEN_2532;
  assign _GEN_2534 = 9'h160 == _T_8348 ? 1'h1 : _GEN_2533;
  assign _GEN_2535 = 9'h161 == _T_8348 ? 1'h1 : _GEN_2534;
  assign _GEN_2536 = 9'h162 == _T_8348 ? 1'h1 : _GEN_2535;
  assign _GEN_2537 = 9'h163 == _T_8348 ? 1'h1 : _GEN_2536;
  assign _GEN_2538 = 9'h164 == _T_8348 ? 1'h1 : _GEN_2537;
  assign _GEN_2539 = 9'h165 == _T_8348 ? 1'h1 : _GEN_2538;
  assign _GEN_2540 = 9'h166 == _T_8348 ? 1'h1 : _GEN_2539;
  assign _GEN_2541 = 9'h167 == _T_8348 ? 1'h1 : _GEN_2540;
  assign _GEN_2542 = 9'h168 == _T_8348 ? 1'h1 : _GEN_2541;
  assign _GEN_2543 = 9'h169 == _T_8348 ? 1'h1 : _GEN_2542;
  assign _GEN_2544 = 9'h16a == _T_8348 ? 1'h1 : _GEN_2543;
  assign _GEN_2545 = 9'h16b == _T_8348 ? 1'h1 : _GEN_2544;
  assign _GEN_2546 = 9'h16c == _T_8348 ? 1'h1 : _GEN_2545;
  assign _GEN_2547 = 9'h16d == _T_8348 ? 1'h1 : _GEN_2546;
  assign _GEN_2548 = 9'h16e == _T_8348 ? 1'h1 : _GEN_2547;
  assign _GEN_2549 = 9'h16f == _T_8348 ? 1'h1 : _GEN_2548;
  assign _GEN_2550 = 9'h170 == _T_8348 ? 1'h1 : _GEN_2549;
  assign _GEN_2551 = 9'h171 == _T_8348 ? 1'h1 : _GEN_2550;
  assign _GEN_2552 = 9'h172 == _T_8348 ? 1'h1 : _GEN_2551;
  assign _GEN_2553 = 9'h173 == _T_8348 ? 1'h1 : _GEN_2552;
  assign _GEN_2554 = 9'h174 == _T_8348 ? 1'h1 : _GEN_2553;
  assign _GEN_2555 = 9'h175 == _T_8348 ? 1'h1 : _GEN_2554;
  assign _GEN_2556 = 9'h176 == _T_8348 ? 1'h1 : _GEN_2555;
  assign _GEN_2557 = 9'h177 == _T_8348 ? 1'h1 : _GEN_2556;
  assign _GEN_2558 = 9'h178 == _T_8348 ? 1'h1 : _GEN_2557;
  assign _GEN_2559 = 9'h179 == _T_8348 ? 1'h1 : _GEN_2558;
  assign _GEN_2560 = 9'h17a == _T_8348 ? 1'h1 : _GEN_2559;
  assign _GEN_2561 = 9'h17b == _T_8348 ? 1'h1 : _GEN_2560;
  assign _GEN_2562 = 9'h17c == _T_8348 ? 1'h1 : _GEN_2561;
  assign _GEN_2563 = 9'h17d == _T_8348 ? 1'h1 : _GEN_2562;
  assign _GEN_2564 = 9'h17e == _T_8348 ? 1'h1 : _GEN_2563;
  assign _GEN_2565 = 9'h17f == _T_8348 ? 1'h1 : _GEN_2564;
  assign _GEN_2566 = 9'h180 == _T_8348 ? 1'h1 : _GEN_2565;
  assign _GEN_2567 = 9'h181 == _T_8348 ? 1'h1 : _GEN_2566;
  assign _GEN_2568 = 9'h182 == _T_8348 ? 1'h1 : _GEN_2567;
  assign _GEN_2569 = 9'h183 == _T_8348 ? 1'h1 : _GEN_2568;
  assign _GEN_2570 = 9'h184 == _T_8348 ? 1'h1 : _GEN_2569;
  assign _GEN_2571 = 9'h185 == _T_8348 ? 1'h1 : _GEN_2570;
  assign _GEN_2572 = 9'h186 == _T_8348 ? 1'h1 : _GEN_2571;
  assign _GEN_2573 = 9'h187 == _T_8348 ? 1'h1 : _GEN_2572;
  assign _GEN_2574 = 9'h188 == _T_8348 ? 1'h1 : _GEN_2573;
  assign _GEN_2575 = 9'h189 == _T_8348 ? 1'h1 : _GEN_2574;
  assign _GEN_2576 = 9'h18a == _T_8348 ? 1'h1 : _GEN_2575;
  assign _GEN_2577 = 9'h18b == _T_8348 ? 1'h1 : _GEN_2576;
  assign _GEN_2578 = 9'h18c == _T_8348 ? 1'h1 : _GEN_2577;
  assign _GEN_2579 = 9'h18d == _T_8348 ? 1'h1 : _GEN_2578;
  assign _GEN_2580 = 9'h18e == _T_8348 ? 1'h1 : _GEN_2579;
  assign _GEN_2581 = 9'h18f == _T_8348 ? 1'h1 : _GEN_2580;
  assign _GEN_2582 = 9'h190 == _T_8348 ? 1'h1 : _GEN_2581;
  assign _GEN_2583 = 9'h191 == _T_8348 ? 1'h1 : _GEN_2582;
  assign _GEN_2584 = 9'h192 == _T_8348 ? 1'h1 : _GEN_2583;
  assign _GEN_2585 = 9'h193 == _T_8348 ? 1'h1 : _GEN_2584;
  assign _GEN_2586 = 9'h194 == _T_8348 ? 1'h1 : _GEN_2585;
  assign _GEN_2587 = 9'h195 == _T_8348 ? 1'h1 : _GEN_2586;
  assign _GEN_2588 = 9'h196 == _T_8348 ? 1'h1 : _GEN_2587;
  assign _GEN_2589 = 9'h197 == _T_8348 ? 1'h1 : _GEN_2588;
  assign _GEN_2590 = 9'h198 == _T_8348 ? 1'h1 : _GEN_2589;
  assign _GEN_2591 = 9'h199 == _T_8348 ? 1'h1 : _GEN_2590;
  assign _GEN_2592 = 9'h19a == _T_8348 ? 1'h1 : _GEN_2591;
  assign _GEN_2593 = 9'h19b == _T_8348 ? 1'h1 : _GEN_2592;
  assign _GEN_2594 = 9'h19c == _T_8348 ? 1'h1 : _GEN_2593;
  assign _GEN_2595 = 9'h19d == _T_8348 ? 1'h1 : _GEN_2594;
  assign _GEN_2596 = 9'h19e == _T_8348 ? 1'h1 : _GEN_2595;
  assign _GEN_2597 = 9'h19f == _T_8348 ? 1'h1 : _GEN_2596;
  assign _GEN_2598 = 9'h1a0 == _T_8348 ? 1'h1 : _GEN_2597;
  assign _GEN_2599 = 9'h1a1 == _T_8348 ? 1'h1 : _GEN_2598;
  assign _GEN_2600 = 9'h1a2 == _T_8348 ? 1'h1 : _GEN_2599;
  assign _GEN_2601 = 9'h1a3 == _T_8348 ? 1'h1 : _GEN_2600;
  assign _GEN_2602 = 9'h1a4 == _T_8348 ? 1'h1 : _GEN_2601;
  assign _GEN_2603 = 9'h1a5 == _T_8348 ? 1'h1 : _GEN_2602;
  assign _GEN_2604 = 9'h1a6 == _T_8348 ? 1'h1 : _GEN_2603;
  assign _GEN_2605 = 9'h1a7 == _T_8348 ? 1'h1 : _GEN_2604;
  assign _GEN_2606 = 9'h1a8 == _T_8348 ? 1'h1 : _GEN_2605;
  assign _GEN_2607 = 9'h1a9 == _T_8348 ? 1'h1 : _GEN_2606;
  assign _GEN_2608 = 9'h1aa == _T_8348 ? 1'h1 : _GEN_2607;
  assign _GEN_2609 = 9'h1ab == _T_8348 ? 1'h1 : _GEN_2608;
  assign _GEN_2610 = 9'h1ac == _T_8348 ? 1'h1 : _GEN_2609;
  assign _GEN_2611 = 9'h1ad == _T_8348 ? 1'h1 : _GEN_2610;
  assign _GEN_2612 = 9'h1ae == _T_8348 ? 1'h1 : _GEN_2611;
  assign _GEN_2613 = 9'h1af == _T_8348 ? 1'h1 : _GEN_2612;
  assign _GEN_2614 = 9'h1b0 == _T_8348 ? 1'h1 : _GEN_2613;
  assign _GEN_2615 = 9'h1b1 == _T_8348 ? 1'h1 : _GEN_2614;
  assign _GEN_2616 = 9'h1b2 == _T_8348 ? 1'h1 : _GEN_2615;
  assign _GEN_2617 = 9'h1b3 == _T_8348 ? 1'h1 : _GEN_2616;
  assign _GEN_2618 = 9'h1b4 == _T_8348 ? 1'h1 : _GEN_2617;
  assign _GEN_2619 = 9'h1b5 == _T_8348 ? 1'h1 : _GEN_2618;
  assign _GEN_2620 = 9'h1b6 == _T_8348 ? 1'h1 : _GEN_2619;
  assign _GEN_2621 = 9'h1b7 == _T_8348 ? 1'h1 : _GEN_2620;
  assign _GEN_2622 = 9'h1b8 == _T_8348 ? 1'h1 : _GEN_2621;
  assign _GEN_2623 = 9'h1b9 == _T_8348 ? 1'h1 : _GEN_2622;
  assign _GEN_2624 = 9'h1ba == _T_8348 ? 1'h1 : _GEN_2623;
  assign _GEN_2625 = 9'h1bb == _T_8348 ? 1'h1 : _GEN_2624;
  assign _GEN_2626 = 9'h1bc == _T_8348 ? 1'h1 : _GEN_2625;
  assign _GEN_2627 = 9'h1bd == _T_8348 ? 1'h1 : _GEN_2626;
  assign _GEN_2628 = 9'h1be == _T_8348 ? 1'h1 : _GEN_2627;
  assign _GEN_2629 = 9'h1bf == _T_8348 ? 1'h1 : _GEN_2628;
  assign _GEN_2630 = 9'h1c0 == _T_8348 ? 1'h1 : _GEN_2629;
  assign _GEN_2631 = 9'h1c1 == _T_8348 ? 1'h1 : _GEN_2630;
  assign _GEN_2632 = 9'h1c2 == _T_8348 ? 1'h1 : _GEN_2631;
  assign _GEN_2633 = 9'h1c3 == _T_8348 ? 1'h1 : _GEN_2632;
  assign _GEN_2634 = 9'h1c4 == _T_8348 ? 1'h1 : _GEN_2633;
  assign _GEN_2635 = 9'h1c5 == _T_8348 ? 1'h1 : _GEN_2634;
  assign _GEN_2636 = 9'h1c6 == _T_8348 ? 1'h1 : _GEN_2635;
  assign _GEN_2637 = 9'h1c7 == _T_8348 ? 1'h1 : _GEN_2636;
  assign _GEN_2638 = 9'h1c8 == _T_8348 ? 1'h1 : _GEN_2637;
  assign _GEN_2639 = 9'h1c9 == _T_8348 ? 1'h1 : _GEN_2638;
  assign _GEN_2640 = 9'h1ca == _T_8348 ? 1'h1 : _GEN_2639;
  assign _GEN_2641 = 9'h1cb == _T_8348 ? 1'h1 : _GEN_2640;
  assign _GEN_2642 = 9'h1cc == _T_8348 ? 1'h1 : _GEN_2641;
  assign _GEN_2643 = 9'h1cd == _T_8348 ? 1'h1 : _GEN_2642;
  assign _GEN_2644 = 9'h1ce == _T_8348 ? 1'h1 : _GEN_2643;
  assign _GEN_2645 = 9'h1cf == _T_8348 ? 1'h1 : _GEN_2644;
  assign _GEN_2646 = 9'h1d0 == _T_8348 ? 1'h1 : _GEN_2645;
  assign _GEN_2647 = 9'h1d1 == _T_8348 ? 1'h1 : _GEN_2646;
  assign _GEN_2648 = 9'h1d2 == _T_8348 ? 1'h1 : _GEN_2647;
  assign _GEN_2649 = 9'h1d3 == _T_8348 ? 1'h1 : _GEN_2648;
  assign _GEN_2650 = 9'h1d4 == _T_8348 ? 1'h1 : _GEN_2649;
  assign _GEN_2651 = 9'h1d5 == _T_8348 ? 1'h1 : _GEN_2650;
  assign _GEN_2652 = 9'h1d6 == _T_8348 ? 1'h1 : _GEN_2651;
  assign _GEN_2653 = 9'h1d7 == _T_8348 ? 1'h1 : _GEN_2652;
  assign _GEN_2654 = 9'h1d8 == _T_8348 ? 1'h1 : _GEN_2653;
  assign _GEN_2655 = 9'h1d9 == _T_8348 ? 1'h1 : _GEN_2654;
  assign _GEN_2656 = 9'h1da == _T_8348 ? 1'h1 : _GEN_2655;
  assign _GEN_2657 = 9'h1db == _T_8348 ? 1'h1 : _GEN_2656;
  assign _GEN_2658 = 9'h1dc == _T_8348 ? 1'h1 : _GEN_2657;
  assign _GEN_2659 = 9'h1dd == _T_8348 ? 1'h1 : _GEN_2658;
  assign _GEN_2660 = 9'h1de == _T_8348 ? 1'h1 : _GEN_2659;
  assign _GEN_2661 = 9'h1df == _T_8348 ? 1'h1 : _GEN_2660;
  assign _GEN_2662 = 9'h1e0 == _T_8348 ? 1'h1 : _GEN_2661;
  assign _GEN_2663 = 9'h1e1 == _T_8348 ? 1'h1 : _GEN_2662;
  assign _GEN_2664 = 9'h1e2 == _T_8348 ? 1'h1 : _GEN_2663;
  assign _GEN_2665 = 9'h1e3 == _T_8348 ? 1'h1 : _GEN_2664;
  assign _GEN_2666 = 9'h1e4 == _T_8348 ? 1'h1 : _GEN_2665;
  assign _GEN_2667 = 9'h1e5 == _T_8348 ? 1'h1 : _GEN_2666;
  assign _GEN_2668 = 9'h1e6 == _T_8348 ? 1'h1 : _GEN_2667;
  assign _GEN_2669 = 9'h1e7 == _T_8348 ? 1'h1 : _GEN_2668;
  assign _GEN_2670 = 9'h1e8 == _T_8348 ? 1'h1 : _GEN_2669;
  assign _GEN_2671 = 9'h1e9 == _T_8348 ? 1'h1 : _GEN_2670;
  assign _GEN_2672 = 9'h1ea == _T_8348 ? 1'h1 : _GEN_2671;
  assign _GEN_2673 = 9'h1eb == _T_8348 ? 1'h1 : _GEN_2672;
  assign _GEN_2674 = 9'h1ec == _T_8348 ? 1'h1 : _GEN_2673;
  assign _GEN_2675 = 9'h1ed == _T_8348 ? 1'h1 : _GEN_2674;
  assign _GEN_2676 = 9'h1ee == _T_8348 ? 1'h1 : _GEN_2675;
  assign _GEN_2677 = 9'h1ef == _T_8348 ? 1'h1 : _GEN_2676;
  assign _GEN_2678 = 9'h1f0 == _T_8348 ? 1'h1 : _GEN_2677;
  assign _GEN_2679 = 9'h1f1 == _T_8348 ? 1'h1 : _GEN_2678;
  assign _GEN_2680 = 9'h1f2 == _T_8348 ? 1'h1 : _GEN_2679;
  assign _GEN_2681 = 9'h1f3 == _T_8348 ? 1'h1 : _GEN_2680;
  assign _GEN_2682 = 9'h1f4 == _T_8348 ? 1'h1 : _GEN_2681;
  assign _GEN_2683 = 9'h1f5 == _T_8348 ? 1'h1 : _GEN_2682;
  assign _GEN_2684 = 9'h1f6 == _T_8348 ? 1'h1 : _GEN_2683;
  assign _GEN_2685 = 9'h1f7 == _T_8348 ? 1'h1 : _GEN_2684;
  assign _GEN_2686 = 9'h1f8 == _T_8348 ? 1'h1 : _GEN_2685;
  assign _GEN_2687 = 9'h1f9 == _T_8348 ? 1'h1 : _GEN_2686;
  assign _GEN_2688 = 9'h1fa == _T_8348 ? 1'h1 : _GEN_2687;
  assign _GEN_2689 = 9'h1fb == _T_8348 ? 1'h1 : _GEN_2688;
  assign _GEN_2690 = 9'h1fc == _T_8348 ? 1'h1 : _GEN_2689;
  assign _GEN_2691 = 9'h1fd == _T_8348 ? 1'h1 : _GEN_2690;
  assign _GEN_2692 = 9'h1fe == _T_8348 ? 1'h1 : _GEN_2691;
  assign _GEN_2693 = 9'h1ff == _T_8348 ? 1'h1 : _GEN_2692;
  assign _GEN_2694 = 9'h1 == _T_8348 ? _T_28371_1 : 32'h0;
  assign _GEN_2695 = 9'h2 == _T_8348 ? _T_28371_2 : _GEN_2694;
  assign _GEN_2696 = 9'h3 == _T_8348 ? _T_28371_3 : _GEN_2695;
  assign _GEN_2697 = 9'h4 == _T_8348 ? _T_28371_4 : _GEN_2696;
  assign _GEN_2698 = 9'h5 == _T_8348 ? _T_28371_5 : _GEN_2697;
  assign _GEN_2699 = 9'h6 == _T_8348 ? _T_28371_6 : _GEN_2698;
  assign _GEN_2700 = 9'h7 == _T_8348 ? _T_28371_7 : _GEN_2699;
  assign _GEN_2701 = 9'h8 == _T_8348 ? _T_28371_8 : _GEN_2700;
  assign _GEN_2702 = 9'h9 == _T_8348 ? _T_28371_9 : _GEN_2701;
  assign _GEN_2703 = 9'ha == _T_8348 ? _T_28371_10 : _GEN_2702;
  assign _GEN_2704 = 9'hb == _T_8348 ? _T_28371_11 : _GEN_2703;
  assign _GEN_2705 = 9'hc == _T_8348 ? _T_28371_12 : _GEN_2704;
  assign _GEN_2706 = 9'hd == _T_8348 ? _T_28371_13 : _GEN_2705;
  assign _GEN_2707 = 9'he == _T_8348 ? _T_28371_14 : _GEN_2706;
  assign _GEN_2708 = 9'hf == _T_8348 ? _T_28371_15 : _GEN_2707;
  assign _GEN_2709 = 9'h10 == _T_8348 ? _T_28371_16 : _GEN_2708;
  assign _GEN_2710 = 9'h11 == _T_8348 ? _T_28371_17 : _GEN_2709;
  assign _GEN_2711 = 9'h12 == _T_8348 ? _T_28371_18 : _GEN_2710;
  assign _GEN_2712 = 9'h13 == _T_8348 ? _T_28371_19 : _GEN_2711;
  assign _GEN_2713 = 9'h14 == _T_8348 ? _T_28371_20 : _GEN_2712;
  assign _GEN_2714 = 9'h15 == _T_8348 ? _T_28371_21 : _GEN_2713;
  assign _GEN_2715 = 9'h16 == _T_8348 ? _T_28371_22 : _GEN_2714;
  assign _GEN_2716 = 9'h17 == _T_8348 ? _T_28371_23 : _GEN_2715;
  assign _GEN_2717 = 9'h18 == _T_8348 ? _T_28371_24 : _GEN_2716;
  assign _GEN_2718 = 9'h19 == _T_8348 ? _T_28371_25 : _GEN_2717;
  assign _GEN_2719 = 9'h1a == _T_8348 ? _T_28371_26 : _GEN_2718;
  assign _GEN_2720 = 9'h1b == _T_8348 ? _T_28371_27 : _GEN_2719;
  assign _GEN_2721 = 9'h1c == _T_8348 ? _T_28371_28 : _GEN_2720;
  assign _GEN_2722 = 9'h1d == _T_8348 ? _T_28371_29 : _GEN_2721;
  assign _GEN_2723 = 9'h1e == _T_8348 ? _T_28371_30 : _GEN_2722;
  assign _GEN_2724 = 9'h1f == _T_8348 ? _T_28371_31 : _GEN_2723;
  assign _GEN_2725 = 9'h20 == _T_8348 ? _T_28371_32 : _GEN_2724;
  assign _GEN_2726 = 9'h21 == _T_8348 ? 32'h0 : _GEN_2725;
  assign _GEN_2727 = 9'h22 == _T_8348 ? 32'h0 : _GEN_2726;
  assign _GEN_2728 = 9'h23 == _T_8348 ? 32'h0 : _GEN_2727;
  assign _GEN_2729 = 9'h24 == _T_8348 ? 32'h0 : _GEN_2728;
  assign _GEN_2730 = 9'h25 == _T_8348 ? 32'h0 : _GEN_2729;
  assign _GEN_2731 = 9'h26 == _T_8348 ? 32'h0 : _GEN_2730;
  assign _GEN_2732 = 9'h27 == _T_8348 ? 32'h0 : _GEN_2731;
  assign _GEN_2733 = 9'h28 == _T_8348 ? 32'h0 : _GEN_2732;
  assign _GEN_2734 = 9'h29 == _T_8348 ? 32'h0 : _GEN_2733;
  assign _GEN_2735 = 9'h2a == _T_8348 ? 32'h0 : _GEN_2734;
  assign _GEN_2736 = 9'h2b == _T_8348 ? 32'h0 : _GEN_2735;
  assign _GEN_2737 = 9'h2c == _T_8348 ? 32'h0 : _GEN_2736;
  assign _GEN_2738 = 9'h2d == _T_8348 ? 32'h0 : _GEN_2737;
  assign _GEN_2739 = 9'h2e == _T_8348 ? 32'h0 : _GEN_2738;
  assign _GEN_2740 = 9'h2f == _T_8348 ? 32'h0 : _GEN_2739;
  assign _GEN_2741 = 9'h30 == _T_8348 ? 32'h0 : _GEN_2740;
  assign _GEN_2742 = 9'h31 == _T_8348 ? 32'h0 : _GEN_2741;
  assign _GEN_2743 = 9'h32 == _T_8348 ? 32'h0 : _GEN_2742;
  assign _GEN_2744 = 9'h33 == _T_8348 ? 32'h0 : _GEN_2743;
  assign _GEN_2745 = 9'h34 == _T_8348 ? 32'h0 : _GEN_2744;
  assign _GEN_2746 = 9'h35 == _T_8348 ? 32'h0 : _GEN_2745;
  assign _GEN_2747 = 9'h36 == _T_8348 ? 32'h0 : _GEN_2746;
  assign _GEN_2748 = 9'h37 == _T_8348 ? 32'h0 : _GEN_2747;
  assign _GEN_2749 = 9'h38 == _T_8348 ? 32'h0 : _GEN_2748;
  assign _GEN_2750 = 9'h39 == _T_8348 ? 32'h0 : _GEN_2749;
  assign _GEN_2751 = 9'h3a == _T_8348 ? 32'h0 : _GEN_2750;
  assign _GEN_2752 = 9'h3b == _T_8348 ? 32'h0 : _GEN_2751;
  assign _GEN_2753 = 9'h3c == _T_8348 ? 32'h0 : _GEN_2752;
  assign _GEN_2754 = 9'h3d == _T_8348 ? 32'h0 : _GEN_2753;
  assign _GEN_2755 = 9'h3e == _T_8348 ? 32'h0 : _GEN_2754;
  assign _GEN_2756 = 9'h3f == _T_8348 ? 32'h0 : _GEN_2755;
  assign _GEN_2757 = 9'h40 == _T_8348 ? _T_28371_64 : _GEN_2756;
  assign _GEN_2758 = 9'h41 == _T_8348 ? _T_28371_65 : _GEN_2757;
  assign _GEN_2759 = 9'h42 == _T_8348 ? 32'h0 : _GEN_2758;
  assign _GEN_2760 = 9'h43 == _T_8348 ? 32'h0 : _GEN_2759;
  assign _GEN_2761 = 9'h44 == _T_8348 ? 32'h0 : _GEN_2760;
  assign _GEN_2762 = 9'h45 == _T_8348 ? 32'h0 : _GEN_2761;
  assign _GEN_2763 = 9'h46 == _T_8348 ? 32'h0 : _GEN_2762;
  assign _GEN_2764 = 9'h47 == _T_8348 ? 32'h0 : _GEN_2763;
  assign _GEN_2765 = 9'h48 == _T_8348 ? 32'h0 : _GEN_2764;
  assign _GEN_2766 = 9'h49 == _T_8348 ? 32'h0 : _GEN_2765;
  assign _GEN_2767 = 9'h4a == _T_8348 ? 32'h0 : _GEN_2766;
  assign _GEN_2768 = 9'h4b == _T_8348 ? 32'h0 : _GEN_2767;
  assign _GEN_2769 = 9'h4c == _T_8348 ? 32'h0 : _GEN_2768;
  assign _GEN_2770 = 9'h4d == _T_8348 ? 32'h0 : _GEN_2769;
  assign _GEN_2771 = 9'h4e == _T_8348 ? 32'h0 : _GEN_2770;
  assign _GEN_2772 = 9'h4f == _T_8348 ? 32'h0 : _GEN_2771;
  assign _GEN_2773 = 9'h50 == _T_8348 ? 32'h0 : _GEN_2772;
  assign _GEN_2774 = 9'h51 == _T_8348 ? 32'h0 : _GEN_2773;
  assign _GEN_2775 = 9'h52 == _T_8348 ? 32'h0 : _GEN_2774;
  assign _GEN_2776 = 9'h53 == _T_8348 ? 32'h0 : _GEN_2775;
  assign _GEN_2777 = 9'h54 == _T_8348 ? 32'h0 : _GEN_2776;
  assign _GEN_2778 = 9'h55 == _T_8348 ? 32'h0 : _GEN_2777;
  assign _GEN_2779 = 9'h56 == _T_8348 ? 32'h0 : _GEN_2778;
  assign _GEN_2780 = 9'h57 == _T_8348 ? 32'h0 : _GEN_2779;
  assign _GEN_2781 = 9'h58 == _T_8348 ? 32'h0 : _GEN_2780;
  assign _GEN_2782 = 9'h59 == _T_8348 ? 32'h0 : _GEN_2781;
  assign _GEN_2783 = 9'h5a == _T_8348 ? 32'h0 : _GEN_2782;
  assign _GEN_2784 = 9'h5b == _T_8348 ? 32'h0 : _GEN_2783;
  assign _GEN_2785 = 9'h5c == _T_8348 ? 32'h0 : _GEN_2784;
  assign _GEN_2786 = 9'h5d == _T_8348 ? 32'h0 : _GEN_2785;
  assign _GEN_2787 = 9'h5e == _T_8348 ? 32'h0 : _GEN_2786;
  assign _GEN_2788 = 9'h5f == _T_8348 ? 32'h0 : _GEN_2787;
  assign _GEN_2789 = 9'h60 == _T_8348 ? 32'h0 : _GEN_2788;
  assign _GEN_2790 = 9'h61 == _T_8348 ? 32'h0 : _GEN_2789;
  assign _GEN_2791 = 9'h62 == _T_8348 ? 32'h0 : _GEN_2790;
  assign _GEN_2792 = 9'h63 == _T_8348 ? 32'h0 : _GEN_2791;
  assign _GEN_2793 = 9'h64 == _T_8348 ? 32'h0 : _GEN_2792;
  assign _GEN_2794 = 9'h65 == _T_8348 ? 32'h0 : _GEN_2793;
  assign _GEN_2795 = 9'h66 == _T_8348 ? 32'h0 : _GEN_2794;
  assign _GEN_2796 = 9'h67 == _T_8348 ? 32'h0 : _GEN_2795;
  assign _GEN_2797 = 9'h68 == _T_8348 ? 32'h0 : _GEN_2796;
  assign _GEN_2798 = 9'h69 == _T_8348 ? 32'h0 : _GEN_2797;
  assign _GEN_2799 = 9'h6a == _T_8348 ? 32'h0 : _GEN_2798;
  assign _GEN_2800 = 9'h6b == _T_8348 ? 32'h0 : _GEN_2799;
  assign _GEN_2801 = 9'h6c == _T_8348 ? 32'h0 : _GEN_2800;
  assign _GEN_2802 = 9'h6d == _T_8348 ? 32'h0 : _GEN_2801;
  assign _GEN_2803 = 9'h6e == _T_8348 ? 32'h0 : _GEN_2802;
  assign _GEN_2804 = 9'h6f == _T_8348 ? 32'h0 : _GEN_2803;
  assign _GEN_2805 = 9'h70 == _T_8348 ? 32'h0 : _GEN_2804;
  assign _GEN_2806 = 9'h71 == _T_8348 ? 32'h0 : _GEN_2805;
  assign _GEN_2807 = 9'h72 == _T_8348 ? 32'h0 : _GEN_2806;
  assign _GEN_2808 = 9'h73 == _T_8348 ? 32'h0 : _GEN_2807;
  assign _GEN_2809 = 9'h74 == _T_8348 ? 32'h0 : _GEN_2808;
  assign _GEN_2810 = 9'h75 == _T_8348 ? 32'h0 : _GEN_2809;
  assign _GEN_2811 = 9'h76 == _T_8348 ? 32'h0 : _GEN_2810;
  assign _GEN_2812 = 9'h77 == _T_8348 ? 32'h0 : _GEN_2811;
  assign _GEN_2813 = 9'h78 == _T_8348 ? 32'h0 : _GEN_2812;
  assign _GEN_2814 = 9'h79 == _T_8348 ? 32'h0 : _GEN_2813;
  assign _GEN_2815 = 9'h7a == _T_8348 ? 32'h0 : _GEN_2814;
  assign _GEN_2816 = 9'h7b == _T_8348 ? 32'h0 : _GEN_2815;
  assign _GEN_2817 = 9'h7c == _T_8348 ? 32'h0 : _GEN_2816;
  assign _GEN_2818 = 9'h7d == _T_8348 ? 32'h0 : _GEN_2817;
  assign _GEN_2819 = 9'h7e == _T_8348 ? 32'h0 : _GEN_2818;
  assign _GEN_2820 = 9'h7f == _T_8348 ? 32'h0 : _GEN_2819;
  assign _GEN_2821 = 9'h80 == _T_8348 ? _T_28371_128 : _GEN_2820;
  assign _GEN_2822 = 9'h81 == _T_8348 ? _T_28371_129 : _GEN_2821;
  assign _GEN_2823 = 9'h82 == _T_8348 ? 32'h0 : _GEN_2822;
  assign _GEN_2824 = 9'h83 == _T_8348 ? 32'h0 : _GEN_2823;
  assign _GEN_2825 = 9'h84 == _T_8348 ? 32'h0 : _GEN_2824;
  assign _GEN_2826 = 9'h85 == _T_8348 ? 32'h0 : _GEN_2825;
  assign _GEN_2827 = 9'h86 == _T_8348 ? 32'h0 : _GEN_2826;
  assign _GEN_2828 = 9'h87 == _T_8348 ? 32'h0 : _GEN_2827;
  assign _GEN_2829 = 9'h88 == _T_8348 ? 32'h0 : _GEN_2828;
  assign _GEN_2830 = 9'h89 == _T_8348 ? 32'h0 : _GEN_2829;
  assign _GEN_2831 = 9'h8a == _T_8348 ? 32'h0 : _GEN_2830;
  assign _GEN_2832 = 9'h8b == _T_8348 ? 32'h0 : _GEN_2831;
  assign _GEN_2833 = 9'h8c == _T_8348 ? 32'h0 : _GEN_2832;
  assign _GEN_2834 = 9'h8d == _T_8348 ? 32'h0 : _GEN_2833;
  assign _GEN_2835 = 9'h8e == _T_8348 ? 32'h0 : _GEN_2834;
  assign _GEN_2836 = 9'h8f == _T_8348 ? 32'h0 : _GEN_2835;
  assign _GEN_2837 = 9'h90 == _T_8348 ? 32'h0 : _GEN_2836;
  assign _GEN_2838 = 9'h91 == _T_8348 ? 32'h0 : _GEN_2837;
  assign _GEN_2839 = 9'h92 == _T_8348 ? 32'h0 : _GEN_2838;
  assign _GEN_2840 = 9'h93 == _T_8348 ? 32'h0 : _GEN_2839;
  assign _GEN_2841 = 9'h94 == _T_8348 ? 32'h0 : _GEN_2840;
  assign _GEN_2842 = 9'h95 == _T_8348 ? 32'h0 : _GEN_2841;
  assign _GEN_2843 = 9'h96 == _T_8348 ? 32'h0 : _GEN_2842;
  assign _GEN_2844 = 9'h97 == _T_8348 ? 32'h0 : _GEN_2843;
  assign _GEN_2845 = 9'h98 == _T_8348 ? 32'h0 : _GEN_2844;
  assign _GEN_2846 = 9'h99 == _T_8348 ? 32'h0 : _GEN_2845;
  assign _GEN_2847 = 9'h9a == _T_8348 ? 32'h0 : _GEN_2846;
  assign _GEN_2848 = 9'h9b == _T_8348 ? 32'h0 : _GEN_2847;
  assign _GEN_2849 = 9'h9c == _T_8348 ? 32'h0 : _GEN_2848;
  assign _GEN_2850 = 9'h9d == _T_8348 ? 32'h0 : _GEN_2849;
  assign _GEN_2851 = 9'h9e == _T_8348 ? 32'h0 : _GEN_2850;
  assign _GEN_2852 = 9'h9f == _T_8348 ? 32'h0 : _GEN_2851;
  assign _GEN_2853 = 9'ha0 == _T_8348 ? 32'h0 : _GEN_2852;
  assign _GEN_2854 = 9'ha1 == _T_8348 ? 32'h0 : _GEN_2853;
  assign _GEN_2855 = 9'ha2 == _T_8348 ? 32'h0 : _GEN_2854;
  assign _GEN_2856 = 9'ha3 == _T_8348 ? 32'h0 : _GEN_2855;
  assign _GEN_2857 = 9'ha4 == _T_8348 ? 32'h0 : _GEN_2856;
  assign _GEN_2858 = 9'ha5 == _T_8348 ? 32'h0 : _GEN_2857;
  assign _GEN_2859 = 9'ha6 == _T_8348 ? 32'h0 : _GEN_2858;
  assign _GEN_2860 = 9'ha7 == _T_8348 ? 32'h0 : _GEN_2859;
  assign _GEN_2861 = 9'ha8 == _T_8348 ? 32'h0 : _GEN_2860;
  assign _GEN_2862 = 9'ha9 == _T_8348 ? 32'h0 : _GEN_2861;
  assign _GEN_2863 = 9'haa == _T_8348 ? 32'h0 : _GEN_2862;
  assign _GEN_2864 = 9'hab == _T_8348 ? 32'h0 : _GEN_2863;
  assign _GEN_2865 = 9'hac == _T_8348 ? 32'h0 : _GEN_2864;
  assign _GEN_2866 = 9'had == _T_8348 ? 32'h0 : _GEN_2865;
  assign _GEN_2867 = 9'hae == _T_8348 ? 32'h0 : _GEN_2866;
  assign _GEN_2868 = 9'haf == _T_8348 ? 32'h0 : _GEN_2867;
  assign _GEN_2869 = 9'hb0 == _T_8348 ? 32'h0 : _GEN_2868;
  assign _GEN_2870 = 9'hb1 == _T_8348 ? 32'h0 : _GEN_2869;
  assign _GEN_2871 = 9'hb2 == _T_8348 ? 32'h0 : _GEN_2870;
  assign _GEN_2872 = 9'hb3 == _T_8348 ? 32'h0 : _GEN_2871;
  assign _GEN_2873 = 9'hb4 == _T_8348 ? 32'h0 : _GEN_2872;
  assign _GEN_2874 = 9'hb5 == _T_8348 ? 32'h0 : _GEN_2873;
  assign _GEN_2875 = 9'hb6 == _T_8348 ? 32'h0 : _GEN_2874;
  assign _GEN_2876 = 9'hb7 == _T_8348 ? 32'h0 : _GEN_2875;
  assign _GEN_2877 = 9'hb8 == _T_8348 ? 32'h0 : _GEN_2876;
  assign _GEN_2878 = 9'hb9 == _T_8348 ? 32'h0 : _GEN_2877;
  assign _GEN_2879 = 9'hba == _T_8348 ? 32'h0 : _GEN_2878;
  assign _GEN_2880 = 9'hbb == _T_8348 ? 32'h0 : _GEN_2879;
  assign _GEN_2881 = 9'hbc == _T_8348 ? 32'h0 : _GEN_2880;
  assign _GEN_2882 = 9'hbd == _T_8348 ? 32'h0 : _GEN_2881;
  assign _GEN_2883 = 9'hbe == _T_8348 ? 32'h0 : _GEN_2882;
  assign _GEN_2884 = 9'hbf == _T_8348 ? 32'h0 : _GEN_2883;
  assign _GEN_2885 = 9'hc0 == _T_8348 ? 32'h0 : _GEN_2884;
  assign _GEN_2886 = 9'hc1 == _T_8348 ? 32'h0 : _GEN_2885;
  assign _GEN_2887 = 9'hc2 == _T_8348 ? 32'h0 : _GEN_2886;
  assign _GEN_2888 = 9'hc3 == _T_8348 ? 32'h0 : _GEN_2887;
  assign _GEN_2889 = 9'hc4 == _T_8348 ? 32'h0 : _GEN_2888;
  assign _GEN_2890 = 9'hc5 == _T_8348 ? 32'h0 : _GEN_2889;
  assign _GEN_2891 = 9'hc6 == _T_8348 ? 32'h0 : _GEN_2890;
  assign _GEN_2892 = 9'hc7 == _T_8348 ? 32'h0 : _GEN_2891;
  assign _GEN_2893 = 9'hc8 == _T_8348 ? 32'h0 : _GEN_2892;
  assign _GEN_2894 = 9'hc9 == _T_8348 ? 32'h0 : _GEN_2893;
  assign _GEN_2895 = 9'hca == _T_8348 ? 32'h0 : _GEN_2894;
  assign _GEN_2896 = 9'hcb == _T_8348 ? 32'h0 : _GEN_2895;
  assign _GEN_2897 = 9'hcc == _T_8348 ? 32'h0 : _GEN_2896;
  assign _GEN_2898 = 9'hcd == _T_8348 ? 32'h0 : _GEN_2897;
  assign _GEN_2899 = 9'hce == _T_8348 ? 32'h0 : _GEN_2898;
  assign _GEN_2900 = 9'hcf == _T_8348 ? 32'h0 : _GEN_2899;
  assign _GEN_2901 = 9'hd0 == _T_8348 ? 32'h0 : _GEN_2900;
  assign _GEN_2902 = 9'hd1 == _T_8348 ? 32'h0 : _GEN_2901;
  assign _GEN_2903 = 9'hd2 == _T_8348 ? 32'h0 : _GEN_2902;
  assign _GEN_2904 = 9'hd3 == _T_8348 ? 32'h0 : _GEN_2903;
  assign _GEN_2905 = 9'hd4 == _T_8348 ? 32'h0 : _GEN_2904;
  assign _GEN_2906 = 9'hd5 == _T_8348 ? 32'h0 : _GEN_2905;
  assign _GEN_2907 = 9'hd6 == _T_8348 ? 32'h0 : _GEN_2906;
  assign _GEN_2908 = 9'hd7 == _T_8348 ? 32'h0 : _GEN_2907;
  assign _GEN_2909 = 9'hd8 == _T_8348 ? 32'h0 : _GEN_2908;
  assign _GEN_2910 = 9'hd9 == _T_8348 ? 32'h0 : _GEN_2909;
  assign _GEN_2911 = 9'hda == _T_8348 ? 32'h0 : _GEN_2910;
  assign _GEN_2912 = 9'hdb == _T_8348 ? 32'h0 : _GEN_2911;
  assign _GEN_2913 = 9'hdc == _T_8348 ? 32'h0 : _GEN_2912;
  assign _GEN_2914 = 9'hdd == _T_8348 ? 32'h0 : _GEN_2913;
  assign _GEN_2915 = 9'hde == _T_8348 ? 32'h0 : _GEN_2914;
  assign _GEN_2916 = 9'hdf == _T_8348 ? 32'h0 : _GEN_2915;
  assign _GEN_2917 = 9'he0 == _T_8348 ? 32'h0 : _GEN_2916;
  assign _GEN_2918 = 9'he1 == _T_8348 ? 32'h0 : _GEN_2917;
  assign _GEN_2919 = 9'he2 == _T_8348 ? 32'h0 : _GEN_2918;
  assign _GEN_2920 = 9'he3 == _T_8348 ? 32'h0 : _GEN_2919;
  assign _GEN_2921 = 9'he4 == _T_8348 ? 32'h0 : _GEN_2920;
  assign _GEN_2922 = 9'he5 == _T_8348 ? 32'h0 : _GEN_2921;
  assign _GEN_2923 = 9'he6 == _T_8348 ? 32'h0 : _GEN_2922;
  assign _GEN_2924 = 9'he7 == _T_8348 ? 32'h0 : _GEN_2923;
  assign _GEN_2925 = 9'he8 == _T_8348 ? 32'h0 : _GEN_2924;
  assign _GEN_2926 = 9'he9 == _T_8348 ? 32'h0 : _GEN_2925;
  assign _GEN_2927 = 9'hea == _T_8348 ? 32'h0 : _GEN_2926;
  assign _GEN_2928 = 9'heb == _T_8348 ? 32'h0 : _GEN_2927;
  assign _GEN_2929 = 9'hec == _T_8348 ? 32'h0 : _GEN_2928;
  assign _GEN_2930 = 9'hed == _T_8348 ? 32'h0 : _GEN_2929;
  assign _GEN_2931 = 9'hee == _T_8348 ? 32'h0 : _GEN_2930;
  assign _GEN_2932 = 9'hef == _T_8348 ? 32'h0 : _GEN_2931;
  assign _GEN_2933 = 9'hf0 == _T_8348 ? 32'h0 : _GEN_2932;
  assign _GEN_2934 = 9'hf1 == _T_8348 ? 32'h0 : _GEN_2933;
  assign _GEN_2935 = 9'hf2 == _T_8348 ? 32'h0 : _GEN_2934;
  assign _GEN_2936 = 9'hf3 == _T_8348 ? 32'h0 : _GEN_2935;
  assign _GEN_2937 = 9'hf4 == _T_8348 ? 32'h0 : _GEN_2936;
  assign _GEN_2938 = 9'hf5 == _T_8348 ? 32'h0 : _GEN_2937;
  assign _GEN_2939 = 9'hf6 == _T_8348 ? 32'h0 : _GEN_2938;
  assign _GEN_2940 = 9'hf7 == _T_8348 ? 32'h0 : _GEN_2939;
  assign _GEN_2941 = 9'hf8 == _T_8348 ? 32'h0 : _GEN_2940;
  assign _GEN_2942 = 9'hf9 == _T_8348 ? 32'h0 : _GEN_2941;
  assign _GEN_2943 = 9'hfa == _T_8348 ? 32'h0 : _GEN_2942;
  assign _GEN_2944 = 9'hfb == _T_8348 ? 32'h0 : _GEN_2943;
  assign _GEN_2945 = 9'hfc == _T_8348 ? 32'h0 : _GEN_2944;
  assign _GEN_2946 = 9'hfd == _T_8348 ? 32'h0 : _GEN_2945;
  assign _GEN_2947 = 9'hfe == _T_8348 ? 32'h0 : _GEN_2946;
  assign _GEN_2948 = 9'hff == _T_8348 ? 32'h0 : _GEN_2947;
  assign _GEN_2949 = 9'h100 == _T_8348 ? _T_28371_256 : _GEN_2948;
  assign _GEN_2950 = 9'h101 == _T_8348 ? _T_28371_257 : _GEN_2949;
  assign _GEN_2951 = 9'h102 == _T_8348 ? 32'h0 : _GEN_2950;
  assign _GEN_2952 = 9'h103 == _T_8348 ? 32'h0 : _GEN_2951;
  assign _GEN_2953 = 9'h104 == _T_8348 ? 32'h0 : _GEN_2952;
  assign _GEN_2954 = 9'h105 == _T_8348 ? 32'h0 : _GEN_2953;
  assign _GEN_2955 = 9'h106 == _T_8348 ? 32'h0 : _GEN_2954;
  assign _GEN_2956 = 9'h107 == _T_8348 ? 32'h0 : _GEN_2955;
  assign _GEN_2957 = 9'h108 == _T_8348 ? 32'h0 : _GEN_2956;
  assign _GEN_2958 = 9'h109 == _T_8348 ? 32'h0 : _GEN_2957;
  assign _GEN_2959 = 9'h10a == _T_8348 ? 32'h0 : _GEN_2958;
  assign _GEN_2960 = 9'h10b == _T_8348 ? 32'h0 : _GEN_2959;
  assign _GEN_2961 = 9'h10c == _T_8348 ? 32'h0 : _GEN_2960;
  assign _GEN_2962 = 9'h10d == _T_8348 ? 32'h0 : _GEN_2961;
  assign _GEN_2963 = 9'h10e == _T_8348 ? 32'h0 : _GEN_2962;
  assign _GEN_2964 = 9'h10f == _T_8348 ? 32'h0 : _GEN_2963;
  assign _GEN_2965 = 9'h110 == _T_8348 ? 32'h0 : _GEN_2964;
  assign _GEN_2966 = 9'h111 == _T_8348 ? 32'h0 : _GEN_2965;
  assign _GEN_2967 = 9'h112 == _T_8348 ? 32'h0 : _GEN_2966;
  assign _GEN_2968 = 9'h113 == _T_8348 ? 32'h0 : _GEN_2967;
  assign _GEN_2969 = 9'h114 == _T_8348 ? 32'h0 : _GEN_2968;
  assign _GEN_2970 = 9'h115 == _T_8348 ? 32'h0 : _GEN_2969;
  assign _GEN_2971 = 9'h116 == _T_8348 ? 32'h0 : _GEN_2970;
  assign _GEN_2972 = 9'h117 == _T_8348 ? 32'h0 : _GEN_2971;
  assign _GEN_2973 = 9'h118 == _T_8348 ? 32'h0 : _GEN_2972;
  assign _GEN_2974 = 9'h119 == _T_8348 ? 32'h0 : _GEN_2973;
  assign _GEN_2975 = 9'h11a == _T_8348 ? 32'h0 : _GEN_2974;
  assign _GEN_2976 = 9'h11b == _T_8348 ? 32'h0 : _GEN_2975;
  assign _GEN_2977 = 9'h11c == _T_8348 ? 32'h0 : _GEN_2976;
  assign _GEN_2978 = 9'h11d == _T_8348 ? 32'h0 : _GEN_2977;
  assign _GEN_2979 = 9'h11e == _T_8348 ? 32'h0 : _GEN_2978;
  assign _GEN_2980 = 9'h11f == _T_8348 ? 32'h0 : _GEN_2979;
  assign _GEN_2981 = 9'h120 == _T_8348 ? 32'h0 : _GEN_2980;
  assign _GEN_2982 = 9'h121 == _T_8348 ? 32'h0 : _GEN_2981;
  assign _GEN_2983 = 9'h122 == _T_8348 ? 32'h0 : _GEN_2982;
  assign _GEN_2984 = 9'h123 == _T_8348 ? 32'h0 : _GEN_2983;
  assign _GEN_2985 = 9'h124 == _T_8348 ? 32'h0 : _GEN_2984;
  assign _GEN_2986 = 9'h125 == _T_8348 ? 32'h0 : _GEN_2985;
  assign _GEN_2987 = 9'h126 == _T_8348 ? 32'h0 : _GEN_2986;
  assign _GEN_2988 = 9'h127 == _T_8348 ? 32'h0 : _GEN_2987;
  assign _GEN_2989 = 9'h128 == _T_8348 ? 32'h0 : _GEN_2988;
  assign _GEN_2990 = 9'h129 == _T_8348 ? 32'h0 : _GEN_2989;
  assign _GEN_2991 = 9'h12a == _T_8348 ? 32'h0 : _GEN_2990;
  assign _GEN_2992 = 9'h12b == _T_8348 ? 32'h0 : _GEN_2991;
  assign _GEN_2993 = 9'h12c == _T_8348 ? 32'h0 : _GEN_2992;
  assign _GEN_2994 = 9'h12d == _T_8348 ? 32'h0 : _GEN_2993;
  assign _GEN_2995 = 9'h12e == _T_8348 ? 32'h0 : _GEN_2994;
  assign _GEN_2996 = 9'h12f == _T_8348 ? 32'h0 : _GEN_2995;
  assign _GEN_2997 = 9'h130 == _T_8348 ? 32'h0 : _GEN_2996;
  assign _GEN_2998 = 9'h131 == _T_8348 ? 32'h0 : _GEN_2997;
  assign _GEN_2999 = 9'h132 == _T_8348 ? 32'h0 : _GEN_2998;
  assign _GEN_3000 = 9'h133 == _T_8348 ? 32'h0 : _GEN_2999;
  assign _GEN_3001 = 9'h134 == _T_8348 ? 32'h0 : _GEN_3000;
  assign _GEN_3002 = 9'h135 == _T_8348 ? 32'h0 : _GEN_3001;
  assign _GEN_3003 = 9'h136 == _T_8348 ? 32'h0 : _GEN_3002;
  assign _GEN_3004 = 9'h137 == _T_8348 ? 32'h0 : _GEN_3003;
  assign _GEN_3005 = 9'h138 == _T_8348 ? 32'h0 : _GEN_3004;
  assign _GEN_3006 = 9'h139 == _T_8348 ? 32'h0 : _GEN_3005;
  assign _GEN_3007 = 9'h13a == _T_8348 ? 32'h0 : _GEN_3006;
  assign _GEN_3008 = 9'h13b == _T_8348 ? 32'h0 : _GEN_3007;
  assign _GEN_3009 = 9'h13c == _T_8348 ? 32'h0 : _GEN_3008;
  assign _GEN_3010 = 9'h13d == _T_8348 ? 32'h0 : _GEN_3009;
  assign _GEN_3011 = 9'h13e == _T_8348 ? 32'h0 : _GEN_3010;
  assign _GEN_3012 = 9'h13f == _T_8348 ? 32'h0 : _GEN_3011;
  assign _GEN_3013 = 9'h140 == _T_8348 ? 32'h0 : _GEN_3012;
  assign _GEN_3014 = 9'h141 == _T_8348 ? 32'h0 : _GEN_3013;
  assign _GEN_3015 = 9'h142 == _T_8348 ? 32'h0 : _GEN_3014;
  assign _GEN_3016 = 9'h143 == _T_8348 ? 32'h0 : _GEN_3015;
  assign _GEN_3017 = 9'h144 == _T_8348 ? 32'h0 : _GEN_3016;
  assign _GEN_3018 = 9'h145 == _T_8348 ? 32'h0 : _GEN_3017;
  assign _GEN_3019 = 9'h146 == _T_8348 ? 32'h0 : _GEN_3018;
  assign _GEN_3020 = 9'h147 == _T_8348 ? 32'h0 : _GEN_3019;
  assign _GEN_3021 = 9'h148 == _T_8348 ? 32'h0 : _GEN_3020;
  assign _GEN_3022 = 9'h149 == _T_8348 ? 32'h0 : _GEN_3021;
  assign _GEN_3023 = 9'h14a == _T_8348 ? 32'h0 : _GEN_3022;
  assign _GEN_3024 = 9'h14b == _T_8348 ? 32'h0 : _GEN_3023;
  assign _GEN_3025 = 9'h14c == _T_8348 ? 32'h0 : _GEN_3024;
  assign _GEN_3026 = 9'h14d == _T_8348 ? 32'h0 : _GEN_3025;
  assign _GEN_3027 = 9'h14e == _T_8348 ? 32'h0 : _GEN_3026;
  assign _GEN_3028 = 9'h14f == _T_8348 ? 32'h0 : _GEN_3027;
  assign _GEN_3029 = 9'h150 == _T_8348 ? 32'h0 : _GEN_3028;
  assign _GEN_3030 = 9'h151 == _T_8348 ? 32'h0 : _GEN_3029;
  assign _GEN_3031 = 9'h152 == _T_8348 ? 32'h0 : _GEN_3030;
  assign _GEN_3032 = 9'h153 == _T_8348 ? 32'h0 : _GEN_3031;
  assign _GEN_3033 = 9'h154 == _T_8348 ? 32'h0 : _GEN_3032;
  assign _GEN_3034 = 9'h155 == _T_8348 ? 32'h0 : _GEN_3033;
  assign _GEN_3035 = 9'h156 == _T_8348 ? 32'h0 : _GEN_3034;
  assign _GEN_3036 = 9'h157 == _T_8348 ? 32'h0 : _GEN_3035;
  assign _GEN_3037 = 9'h158 == _T_8348 ? 32'h0 : _GEN_3036;
  assign _GEN_3038 = 9'h159 == _T_8348 ? 32'h0 : _GEN_3037;
  assign _GEN_3039 = 9'h15a == _T_8348 ? 32'h0 : _GEN_3038;
  assign _GEN_3040 = 9'h15b == _T_8348 ? 32'h0 : _GEN_3039;
  assign _GEN_3041 = 9'h15c == _T_8348 ? 32'h0 : _GEN_3040;
  assign _GEN_3042 = 9'h15d == _T_8348 ? 32'h0 : _GEN_3041;
  assign _GEN_3043 = 9'h15e == _T_8348 ? 32'h0 : _GEN_3042;
  assign _GEN_3044 = 9'h15f == _T_8348 ? 32'h0 : _GEN_3043;
  assign _GEN_3045 = 9'h160 == _T_8348 ? 32'h0 : _GEN_3044;
  assign _GEN_3046 = 9'h161 == _T_8348 ? 32'h0 : _GEN_3045;
  assign _GEN_3047 = 9'h162 == _T_8348 ? 32'h0 : _GEN_3046;
  assign _GEN_3048 = 9'h163 == _T_8348 ? 32'h0 : _GEN_3047;
  assign _GEN_3049 = 9'h164 == _T_8348 ? 32'h0 : _GEN_3048;
  assign _GEN_3050 = 9'h165 == _T_8348 ? 32'h0 : _GEN_3049;
  assign _GEN_3051 = 9'h166 == _T_8348 ? 32'h0 : _GEN_3050;
  assign _GEN_3052 = 9'h167 == _T_8348 ? 32'h0 : _GEN_3051;
  assign _GEN_3053 = 9'h168 == _T_8348 ? 32'h0 : _GEN_3052;
  assign _GEN_3054 = 9'h169 == _T_8348 ? 32'h0 : _GEN_3053;
  assign _GEN_3055 = 9'h16a == _T_8348 ? 32'h0 : _GEN_3054;
  assign _GEN_3056 = 9'h16b == _T_8348 ? 32'h0 : _GEN_3055;
  assign _GEN_3057 = 9'h16c == _T_8348 ? 32'h0 : _GEN_3056;
  assign _GEN_3058 = 9'h16d == _T_8348 ? 32'h0 : _GEN_3057;
  assign _GEN_3059 = 9'h16e == _T_8348 ? 32'h0 : _GEN_3058;
  assign _GEN_3060 = 9'h16f == _T_8348 ? 32'h0 : _GEN_3059;
  assign _GEN_3061 = 9'h170 == _T_8348 ? 32'h0 : _GEN_3060;
  assign _GEN_3062 = 9'h171 == _T_8348 ? 32'h0 : _GEN_3061;
  assign _GEN_3063 = 9'h172 == _T_8348 ? 32'h0 : _GEN_3062;
  assign _GEN_3064 = 9'h173 == _T_8348 ? 32'h0 : _GEN_3063;
  assign _GEN_3065 = 9'h174 == _T_8348 ? 32'h0 : _GEN_3064;
  assign _GEN_3066 = 9'h175 == _T_8348 ? 32'h0 : _GEN_3065;
  assign _GEN_3067 = 9'h176 == _T_8348 ? 32'h0 : _GEN_3066;
  assign _GEN_3068 = 9'h177 == _T_8348 ? 32'h0 : _GEN_3067;
  assign _GEN_3069 = 9'h178 == _T_8348 ? 32'h0 : _GEN_3068;
  assign _GEN_3070 = 9'h179 == _T_8348 ? 32'h0 : _GEN_3069;
  assign _GEN_3071 = 9'h17a == _T_8348 ? 32'h0 : _GEN_3070;
  assign _GEN_3072 = 9'h17b == _T_8348 ? 32'h0 : _GEN_3071;
  assign _GEN_3073 = 9'h17c == _T_8348 ? 32'h0 : _GEN_3072;
  assign _GEN_3074 = 9'h17d == _T_8348 ? 32'h0 : _GEN_3073;
  assign _GEN_3075 = 9'h17e == _T_8348 ? 32'h0 : _GEN_3074;
  assign _GEN_3076 = 9'h17f == _T_8348 ? 32'h0 : _GEN_3075;
  assign _GEN_3077 = 9'h180 == _T_8348 ? 32'h0 : _GEN_3076;
  assign _GEN_3078 = 9'h181 == _T_8348 ? 32'h0 : _GEN_3077;
  assign _GEN_3079 = 9'h182 == _T_8348 ? 32'h0 : _GEN_3078;
  assign _GEN_3080 = 9'h183 == _T_8348 ? 32'h0 : _GEN_3079;
  assign _GEN_3081 = 9'h184 == _T_8348 ? 32'h0 : _GEN_3080;
  assign _GEN_3082 = 9'h185 == _T_8348 ? 32'h0 : _GEN_3081;
  assign _GEN_3083 = 9'h186 == _T_8348 ? 32'h0 : _GEN_3082;
  assign _GEN_3084 = 9'h187 == _T_8348 ? 32'h0 : _GEN_3083;
  assign _GEN_3085 = 9'h188 == _T_8348 ? 32'h0 : _GEN_3084;
  assign _GEN_3086 = 9'h189 == _T_8348 ? 32'h0 : _GEN_3085;
  assign _GEN_3087 = 9'h18a == _T_8348 ? 32'h0 : _GEN_3086;
  assign _GEN_3088 = 9'h18b == _T_8348 ? 32'h0 : _GEN_3087;
  assign _GEN_3089 = 9'h18c == _T_8348 ? 32'h0 : _GEN_3088;
  assign _GEN_3090 = 9'h18d == _T_8348 ? 32'h0 : _GEN_3089;
  assign _GEN_3091 = 9'h18e == _T_8348 ? 32'h0 : _GEN_3090;
  assign _GEN_3092 = 9'h18f == _T_8348 ? 32'h0 : _GEN_3091;
  assign _GEN_3093 = 9'h190 == _T_8348 ? 32'h0 : _GEN_3092;
  assign _GEN_3094 = 9'h191 == _T_8348 ? 32'h0 : _GEN_3093;
  assign _GEN_3095 = 9'h192 == _T_8348 ? 32'h0 : _GEN_3094;
  assign _GEN_3096 = 9'h193 == _T_8348 ? 32'h0 : _GEN_3095;
  assign _GEN_3097 = 9'h194 == _T_8348 ? 32'h0 : _GEN_3096;
  assign _GEN_3098 = 9'h195 == _T_8348 ? 32'h0 : _GEN_3097;
  assign _GEN_3099 = 9'h196 == _T_8348 ? 32'h0 : _GEN_3098;
  assign _GEN_3100 = 9'h197 == _T_8348 ? 32'h0 : _GEN_3099;
  assign _GEN_3101 = 9'h198 == _T_8348 ? 32'h0 : _GEN_3100;
  assign _GEN_3102 = 9'h199 == _T_8348 ? 32'h0 : _GEN_3101;
  assign _GEN_3103 = 9'h19a == _T_8348 ? 32'h0 : _GEN_3102;
  assign _GEN_3104 = 9'h19b == _T_8348 ? 32'h0 : _GEN_3103;
  assign _GEN_3105 = 9'h19c == _T_8348 ? 32'h0 : _GEN_3104;
  assign _GEN_3106 = 9'h19d == _T_8348 ? 32'h0 : _GEN_3105;
  assign _GEN_3107 = 9'h19e == _T_8348 ? 32'h0 : _GEN_3106;
  assign _GEN_3108 = 9'h19f == _T_8348 ? 32'h0 : _GEN_3107;
  assign _GEN_3109 = 9'h1a0 == _T_8348 ? 32'h0 : _GEN_3108;
  assign _GEN_3110 = 9'h1a1 == _T_8348 ? 32'h0 : _GEN_3109;
  assign _GEN_3111 = 9'h1a2 == _T_8348 ? 32'h0 : _GEN_3110;
  assign _GEN_3112 = 9'h1a3 == _T_8348 ? 32'h0 : _GEN_3111;
  assign _GEN_3113 = 9'h1a4 == _T_8348 ? 32'h0 : _GEN_3112;
  assign _GEN_3114 = 9'h1a5 == _T_8348 ? 32'h0 : _GEN_3113;
  assign _GEN_3115 = 9'h1a6 == _T_8348 ? 32'h0 : _GEN_3114;
  assign _GEN_3116 = 9'h1a7 == _T_8348 ? 32'h0 : _GEN_3115;
  assign _GEN_3117 = 9'h1a8 == _T_8348 ? 32'h0 : _GEN_3116;
  assign _GEN_3118 = 9'h1a9 == _T_8348 ? 32'h0 : _GEN_3117;
  assign _GEN_3119 = 9'h1aa == _T_8348 ? 32'h0 : _GEN_3118;
  assign _GEN_3120 = 9'h1ab == _T_8348 ? 32'h0 : _GEN_3119;
  assign _GEN_3121 = 9'h1ac == _T_8348 ? 32'h0 : _GEN_3120;
  assign _GEN_3122 = 9'h1ad == _T_8348 ? 32'h0 : _GEN_3121;
  assign _GEN_3123 = 9'h1ae == _T_8348 ? 32'h0 : _GEN_3122;
  assign _GEN_3124 = 9'h1af == _T_8348 ? 32'h0 : _GEN_3123;
  assign _GEN_3125 = 9'h1b0 == _T_8348 ? 32'h0 : _GEN_3124;
  assign _GEN_3126 = 9'h1b1 == _T_8348 ? 32'h0 : _GEN_3125;
  assign _GEN_3127 = 9'h1b2 == _T_8348 ? 32'h0 : _GEN_3126;
  assign _GEN_3128 = 9'h1b3 == _T_8348 ? 32'h0 : _GEN_3127;
  assign _GEN_3129 = 9'h1b4 == _T_8348 ? 32'h0 : _GEN_3128;
  assign _GEN_3130 = 9'h1b5 == _T_8348 ? 32'h0 : _GEN_3129;
  assign _GEN_3131 = 9'h1b6 == _T_8348 ? 32'h0 : _GEN_3130;
  assign _GEN_3132 = 9'h1b7 == _T_8348 ? 32'h0 : _GEN_3131;
  assign _GEN_3133 = 9'h1b8 == _T_8348 ? 32'h0 : _GEN_3132;
  assign _GEN_3134 = 9'h1b9 == _T_8348 ? 32'h0 : _GEN_3133;
  assign _GEN_3135 = 9'h1ba == _T_8348 ? 32'h0 : _GEN_3134;
  assign _GEN_3136 = 9'h1bb == _T_8348 ? 32'h0 : _GEN_3135;
  assign _GEN_3137 = 9'h1bc == _T_8348 ? 32'h0 : _GEN_3136;
  assign _GEN_3138 = 9'h1bd == _T_8348 ? 32'h0 : _GEN_3137;
  assign _GEN_3139 = 9'h1be == _T_8348 ? 32'h0 : _GEN_3138;
  assign _GEN_3140 = 9'h1bf == _T_8348 ? 32'h0 : _GEN_3139;
  assign _GEN_3141 = 9'h1c0 == _T_8348 ? 32'h0 : _GEN_3140;
  assign _GEN_3142 = 9'h1c1 == _T_8348 ? 32'h0 : _GEN_3141;
  assign _GEN_3143 = 9'h1c2 == _T_8348 ? 32'h0 : _GEN_3142;
  assign _GEN_3144 = 9'h1c3 == _T_8348 ? 32'h0 : _GEN_3143;
  assign _GEN_3145 = 9'h1c4 == _T_8348 ? 32'h0 : _GEN_3144;
  assign _GEN_3146 = 9'h1c5 == _T_8348 ? 32'h0 : _GEN_3145;
  assign _GEN_3147 = 9'h1c6 == _T_8348 ? 32'h0 : _GEN_3146;
  assign _GEN_3148 = 9'h1c7 == _T_8348 ? 32'h0 : _GEN_3147;
  assign _GEN_3149 = 9'h1c8 == _T_8348 ? 32'h0 : _GEN_3148;
  assign _GEN_3150 = 9'h1c9 == _T_8348 ? 32'h0 : _GEN_3149;
  assign _GEN_3151 = 9'h1ca == _T_8348 ? 32'h0 : _GEN_3150;
  assign _GEN_3152 = 9'h1cb == _T_8348 ? 32'h0 : _GEN_3151;
  assign _GEN_3153 = 9'h1cc == _T_8348 ? 32'h0 : _GEN_3152;
  assign _GEN_3154 = 9'h1cd == _T_8348 ? 32'h0 : _GEN_3153;
  assign _GEN_3155 = 9'h1ce == _T_8348 ? 32'h0 : _GEN_3154;
  assign _GEN_3156 = 9'h1cf == _T_8348 ? 32'h0 : _GEN_3155;
  assign _GEN_3157 = 9'h1d0 == _T_8348 ? 32'h0 : _GEN_3156;
  assign _GEN_3158 = 9'h1d1 == _T_8348 ? 32'h0 : _GEN_3157;
  assign _GEN_3159 = 9'h1d2 == _T_8348 ? 32'h0 : _GEN_3158;
  assign _GEN_3160 = 9'h1d3 == _T_8348 ? 32'h0 : _GEN_3159;
  assign _GEN_3161 = 9'h1d4 == _T_8348 ? 32'h0 : _GEN_3160;
  assign _GEN_3162 = 9'h1d5 == _T_8348 ? 32'h0 : _GEN_3161;
  assign _GEN_3163 = 9'h1d6 == _T_8348 ? 32'h0 : _GEN_3162;
  assign _GEN_3164 = 9'h1d7 == _T_8348 ? 32'h0 : _GEN_3163;
  assign _GEN_3165 = 9'h1d8 == _T_8348 ? 32'h0 : _GEN_3164;
  assign _GEN_3166 = 9'h1d9 == _T_8348 ? 32'h0 : _GEN_3165;
  assign _GEN_3167 = 9'h1da == _T_8348 ? 32'h0 : _GEN_3166;
  assign _GEN_3168 = 9'h1db == _T_8348 ? 32'h0 : _GEN_3167;
  assign _GEN_3169 = 9'h1dc == _T_8348 ? 32'h0 : _GEN_3168;
  assign _GEN_3170 = 9'h1dd == _T_8348 ? 32'h0 : _GEN_3169;
  assign _GEN_3171 = 9'h1de == _T_8348 ? 32'h0 : _GEN_3170;
  assign _GEN_3172 = 9'h1df == _T_8348 ? 32'h0 : _GEN_3171;
  assign _GEN_3173 = 9'h1e0 == _T_8348 ? 32'h0 : _GEN_3172;
  assign _GEN_3174 = 9'h1e1 == _T_8348 ? 32'h0 : _GEN_3173;
  assign _GEN_3175 = 9'h1e2 == _T_8348 ? 32'h0 : _GEN_3174;
  assign _GEN_3176 = 9'h1e3 == _T_8348 ? 32'h0 : _GEN_3175;
  assign _GEN_3177 = 9'h1e4 == _T_8348 ? 32'h0 : _GEN_3176;
  assign _GEN_3178 = 9'h1e5 == _T_8348 ? 32'h0 : _GEN_3177;
  assign _GEN_3179 = 9'h1e6 == _T_8348 ? 32'h0 : _GEN_3178;
  assign _GEN_3180 = 9'h1e7 == _T_8348 ? 32'h0 : _GEN_3179;
  assign _GEN_3181 = 9'h1e8 == _T_8348 ? 32'h0 : _GEN_3180;
  assign _GEN_3182 = 9'h1e9 == _T_8348 ? 32'h0 : _GEN_3181;
  assign _GEN_3183 = 9'h1ea == _T_8348 ? 32'h0 : _GEN_3182;
  assign _GEN_3184 = 9'h1eb == _T_8348 ? 32'h0 : _GEN_3183;
  assign _GEN_3185 = 9'h1ec == _T_8348 ? 32'h0 : _GEN_3184;
  assign _GEN_3186 = 9'h1ed == _T_8348 ? 32'h0 : _GEN_3185;
  assign _GEN_3187 = 9'h1ee == _T_8348 ? 32'h0 : _GEN_3186;
  assign _GEN_3188 = 9'h1ef == _T_8348 ? 32'h0 : _GEN_3187;
  assign _GEN_3189 = 9'h1f0 == _T_8348 ? 32'h0 : _GEN_3188;
  assign _GEN_3190 = 9'h1f1 == _T_8348 ? 32'h0 : _GEN_3189;
  assign _GEN_3191 = 9'h1f2 == _T_8348 ? 32'h0 : _GEN_3190;
  assign _GEN_3192 = 9'h1f3 == _T_8348 ? 32'h0 : _GEN_3191;
  assign _GEN_3193 = 9'h1f4 == _T_8348 ? 32'h0 : _GEN_3192;
  assign _GEN_3194 = 9'h1f5 == _T_8348 ? 32'h0 : _GEN_3193;
  assign _GEN_3195 = 9'h1f6 == _T_8348 ? 32'h0 : _GEN_3194;
  assign _GEN_3196 = 9'h1f7 == _T_8348 ? 32'h0 : _GEN_3195;
  assign _GEN_3197 = 9'h1f8 == _T_8348 ? 32'h0 : _GEN_3196;
  assign _GEN_3198 = 9'h1f9 == _T_8348 ? 32'h0 : _GEN_3197;
  assign _GEN_3199 = 9'h1fa == _T_8348 ? 32'h0 : _GEN_3198;
  assign _GEN_3200 = 9'h1fb == _T_8348 ? 32'h0 : _GEN_3199;
  assign _GEN_3201 = 9'h1fc == _T_8348 ? 32'h0 : _GEN_3200;
  assign _GEN_3202 = 9'h1fd == _T_8348 ? 32'h0 : _GEN_3201;
  assign _GEN_3203 = 9'h1fe == _T_8348 ? 32'h0 : _GEN_3202;
  assign _GEN_3204 = 9'h1ff == _T_8348 ? 32'h0 : _GEN_3203;
  assign _T_28888 = _GEN_5 ? _GEN_6 : 32'h0;
  assign _T_28889 = _T_1859_bits_extra[11:2];
  assign _T_28890 = _T_1859_bits_extra[1:0];
  assign rvx_port_22 = rvx_signal_448;
  assign rvx_port_40 = _T_31_a_ready;
  assign rvx_port_27 = _T_31_d_valid;
  assign rvx_port_39 = _T_31_d_bits_opcode;
  assign rvx_port_14 = _T_31_d_bits_size;
  assign rvx_port_46 = _T_31_d_bits_source;
  assign rvx_port_24 = _T_31_d_bits_data;
  assign _T_31_a_ready = _T_1846_ready;
  assign _T_31_a_valid = rvx_port_34;
  assign _T_31_a_bits_opcode = rvx_port_18;
  assign _T_31_a_bits_size = rvx_port_04;
  assign _T_31_a_bits_source = rvx_port_42;
  assign _T_31_a_bits_address = rvx_port_45;
  assign _T_31_a_bits_mask = rvx_port_38;
  assign _T_31_a_bits_data = rvx_port_33;
  assign _T_31_d_ready = rvx_port_31;
  assign _T_31_d_valid = _T_1859_valid;
  assign _T_31_d_bits_opcode = {{2'd0}, _T_1859_bits_read};
  assign _T_31_d_bits_size = _T_28893_size;
  assign _T_31_d_bits_source = _T_28893_source;
  assign _T_31_d_bits_data = _T_1859_bits_data;
  assign rvx_signal_455 = rvx_port_26;
  assign rvx_signal_394 = rvx_port_03;
  assign rvx_signal_082 = rvx_port_30;
  assign rvx_signal_031 = rvx_port_35;
  assign rvx_signal_112 = rvx_port_13;
  assign rvx_signal_169 = rvx_port_19;
  assign rvx_signal_288 = rvx_port_29;
  assign rvx_signal_353 = rvx_port_32;
  assign rvx_signal_216 = rvx_port_28;
  assign rvx_signal_419 = rvx_port_17;
  assign rvx_signal_109 = rvx_port_12;
  assign rvx_signal_458 = rvx_port_48;
  assign rvx_signal_411 = rvx_port_37;
  assign rvx_signal_412 = rvx_port_43;
  assign rvx_signal_262 = rvx_port_01;
  assign rvx_signal_367 = rvx_port_09;
  assign rvx_signal_200 = rvx_port_05;
  assign rvx_signal_046 = rvx_port_08;
  assign rvx_signal_403 = rvx_port_11;
  assign rvx_signal_402 = rvx_port_47;
  assign rvx_signal_193 = rvx_port_15;
  assign rvx_signal_154 = rvx_port_07;
  assign rvx_signal_325 = rvx_port_23;
  assign rvx_signal_381 = rvx_port_36;
  assign rvx_signal_348 = rvx_port_10;
  assign rvx_signal_334 = rvx_port_06;
  assign rvx_signal_102 = rvx_port_20;
  assign rvx_signal_323 = rvx_port_44;
  assign rvx_signal_231 = rvx_port_02;
  assign rvx_signal_115 = rvx_port_00;
  assign rvx_signal_218 = rvx_port_21;
  assign rvx_signal_122 = rvx_port_16;
  assign rvx_signal_448 = _T_1520;
  assign rvx_signal_123 = 1'h0;
  assign rvx_signal_256 = 1'h1;
  assign rvx_signal_130 = rvx_signal_280;
  assign rvx_signal_108 = rvx_port_25;
  assign rvx_signal_006 = rvx_port_41;
  assign rvx_signal_149 = rvx_signal_455;
  assign rvx_signal_075 = rvx_signal_047;
  assign rvx_signal_027 = rvx_signal_158;
  assign rvx_signal_098 = rvx_port_25;
  assign rvx_signal_081 = rvx_port_41;
  assign rvx_signal_441 = rvx_signal_394;
  assign rvx_signal_452 = rvx_signal_414;
  assign rvx_signal_428 = rvx_signal_357;
  assign rvx_signal_012 = rvx_port_25;
  assign rvx_signal_327 = rvx_port_41;
  assign rvx_signal_461 = rvx_signal_082;
  assign rvx_signal_101 = rvx_signal_313;
  assign rvx_signal_244 = rvx_signal_055;
  assign rvx_signal_338 = rvx_port_25;
  assign rvx_signal_203 = rvx_port_41;
  assign rvx_signal_000 = rvx_signal_031;
  assign rvx_signal_024 = rvx_signal_170;
  assign rvx_signal_174 = rvx_signal_420;
  assign rvx_signal_159 = rvx_port_25;
  assign rvx_signal_054 = rvx_port_41;
  assign rvx_signal_036 = rvx_signal_112;
  assign rvx_signal_341 = rvx_signal_277;
  assign rvx_signal_209 = rvx_signal_453;
  assign rvx_signal_360 = rvx_port_25;
  assign rvx_signal_297 = rvx_port_41;
  assign rvx_signal_198 = rvx_signal_169;
  assign rvx_signal_326 = rvx_signal_040;
  assign rvx_signal_201 = rvx_signal_377;
  assign rvx_signal_401 = rvx_port_25;
  assign rvx_signal_425 = rvx_port_41;
  assign rvx_signal_063 = rvx_signal_288;
  assign rvx_signal_186 = rvx_signal_447;
  assign rvx_signal_379 = rvx_signal_106;
  assign rvx_signal_451 = rvx_port_25;
  assign rvx_signal_074 = rvx_port_41;
  assign rvx_signal_192 = rvx_signal_353;
  assign rvx_signal_312 = rvx_signal_078;
  assign rvx_signal_282 = rvx_signal_134;
  assign rvx_signal_204 = rvx_port_25;
  assign rvx_signal_405 = rvx_port_41;
  assign rvx_signal_148 = rvx_signal_216;
  assign rvx_signal_180 = rvx_signal_457;
  assign rvx_signal_295 = rvx_signal_138;
  assign rvx_signal_125 = rvx_port_25;
  assign rvx_signal_330 = rvx_port_41;
  assign rvx_signal_336 = rvx_signal_419;
  assign rvx_signal_254 = rvx_signal_472;
  assign rvx_signal_391 = rvx_signal_387;
  assign rvx_signal_085 = rvx_port_25;
  assign rvx_signal_163 = rvx_port_41;
  assign rvx_signal_028 = rvx_signal_109;
  assign rvx_signal_062 = rvx_signal_212;
  assign rvx_signal_220 = rvx_signal_069;
  assign rvx_signal_390 = rvx_port_25;
  assign rvx_signal_439 = rvx_port_41;
  assign rvx_signal_141 = rvx_signal_458;
  assign rvx_signal_226 = rvx_signal_473;
  assign rvx_signal_347 = rvx_signal_160;
  assign rvx_signal_299 = rvx_port_25;
  assign rvx_signal_128 = rvx_port_41;
  assign rvx_signal_213 = rvx_signal_411;
  assign rvx_signal_090 = rvx_signal_397;
  assign rvx_signal_151 = rvx_signal_035;
  assign rvx_signal_070 = rvx_port_25;
  assign rvx_signal_039 = rvx_port_41;
  assign rvx_signal_135 = rvx_signal_412;
  assign rvx_signal_127 = rvx_signal_340;
  assign rvx_signal_206 = rvx_signal_421;
  assign rvx_signal_042 = rvx_port_25;
  assign rvx_signal_464 = rvx_port_41;
  assign rvx_signal_010 = rvx_signal_262;
  assign rvx_signal_053 = rvx_signal_247;
  assign rvx_signal_252 = rvx_signal_333;
  assign rvx_signal_235 = rvx_port_25;
  assign rvx_signal_156 = rvx_port_41;
  assign rvx_signal_227 = rvx_signal_367;
  assign rvx_signal_373 = rvx_signal_274;
  assign rvx_signal_041 = rvx_signal_020;
  assign rvx_signal_044 = rvx_port_25;
  assign rvx_signal_398 = rvx_port_41;
  assign rvx_signal_368 = rvx_signal_200;
  assign rvx_signal_037 = rvx_signal_211;
  assign rvx_signal_356 = rvx_signal_207;
  assign rvx_signal_308 = rvx_port_25;
  assign rvx_signal_463 = rvx_port_41;
  assign rvx_signal_236 = rvx_signal_046;
  assign rvx_signal_093 = rvx_signal_171;
  assign rvx_signal_471 = rvx_signal_354;
  assign rvx_signal_187 = rvx_port_25;
  assign rvx_signal_317 = rvx_port_41;
  assign rvx_signal_301 = rvx_signal_403;
  assign rvx_signal_177 = rvx_signal_071;
  assign rvx_signal_324 = rvx_signal_392;
  assign rvx_signal_413 = rvx_port_25;
  assign rvx_signal_013 = rvx_port_41;
  assign rvx_signal_343 = rvx_signal_402;
  assign rvx_signal_389 = rvx_signal_094;
  assign rvx_signal_337 = rvx_signal_176;
  assign rvx_signal_474 = rvx_port_25;
  assign rvx_signal_107 = rvx_port_41;
  assign rvx_signal_477 = rvx_signal_193;
  assign rvx_signal_030 = rvx_signal_139;
  assign rvx_signal_459 = rvx_signal_264;
  assign rvx_signal_015 = rvx_port_25;
  assign rvx_signal_095 = rvx_port_41;
  assign rvx_signal_194 = rvx_signal_154;
  assign rvx_signal_424 = rvx_signal_191;
  assign rvx_signal_329 = rvx_signal_302;
  assign rvx_signal_468 = rvx_port_25;
  assign rvx_signal_084 = rvx_port_41;
  assign rvx_signal_175 = rvx_signal_325;
  assign rvx_signal_223 = rvx_signal_147;
  assign rvx_signal_205 = rvx_signal_342;
  assign rvx_signal_291 = rvx_port_25;
  assign rvx_signal_051 = rvx_port_41;
  assign rvx_signal_352 = rvx_signal_381;
  assign rvx_signal_442 = rvx_signal_105;
  assign rvx_signal_335 = rvx_signal_467;
  assign rvx_signal_257 = rvx_port_25;
  assign rvx_signal_361 = rvx_port_41;
  assign rvx_signal_438 = rvx_signal_348;
  assign rvx_signal_104 = rvx_signal_396;
  assign rvx_signal_219 = rvx_signal_250;
  assign rvx_signal_417 = rvx_port_25;
  assign rvx_signal_217 = rvx_port_41;
  assign rvx_signal_380 = rvx_signal_334;
  assign rvx_signal_113 = rvx_signal_059;
  assign rvx_signal_310 = rvx_signal_476;
  assign rvx_signal_133 = rvx_port_25;
  assign rvx_signal_142 = rvx_port_41;
  assign rvx_signal_091 = rvx_signal_102;
  assign rvx_signal_346 = rvx_signal_319;
  assign rvx_signal_246 = rvx_signal_026;
  assign rvx_signal_079 = rvx_port_25;
  assign rvx_signal_049 = rvx_port_41;
  assign rvx_signal_355 = rvx_signal_323;
  assign rvx_signal_440 = rvx_signal_260;
  assign rvx_signal_157 = rvx_signal_478;
  assign rvx_signal_214 = rvx_port_25;
  assign rvx_signal_261 = rvx_port_41;
  assign rvx_signal_021 = rvx_signal_231;
  assign rvx_signal_320 = rvx_signal_322;
  assign rvx_signal_076 = rvx_signal_230;
  assign rvx_signal_434 = rvx_port_25;
  assign rvx_signal_293 = rvx_port_41;
  assign rvx_signal_393 = rvx_signal_115;
  assign rvx_signal_270 = rvx_signal_456;
  assign rvx_signal_376 = rvx_signal_232;
  assign rvx_signal_016 = rvx_port_25;
  assign rvx_signal_281 = rvx_port_41;
  assign rvx_signal_121 = rvx_signal_218;
  assign rvx_signal_009 = rvx_signal_061;
  assign rvx_signal_237 = rvx_signal_370;
  assign rvx_signal_375 = rvx_port_25;
  assign rvx_signal_362 = rvx_port_41;
  assign rvx_signal_210 = rvx_signal_122;
  assign rvx_signal_284 = rvx_signal_286;
  assign rvx_signal_073 = rvx_signal_339;
  assign rvx_signal_385 = rvx_port_25;
  assign rvx_signal_331 = rvx_port_41;
  assign rvx_signal_280 = _T_1808;
  assign rvx_signal_269 = rvx_signal_307;
  assign rvx_signal_047 = _T_1626;
  assign rvx_signal_158 = _T_1809;
  assign rvx_signal_119 = rvx_signal_146;
  assign rvx_signal_414 = _T_1631;
  assign rvx_signal_357 = _T_1810;
  assign rvx_signal_184 = rvx_signal_152;
  assign rvx_signal_313 = _T_1636;
  assign rvx_signal_055 = _T_1811;
  assign rvx_signal_251 = rvx_signal_321;
  assign rvx_signal_170 = _T_1641;
  assign rvx_signal_420 = _T_1812;
  assign rvx_signal_199 = rvx_signal_100;
  assign rvx_signal_277 = _T_1646;
  assign rvx_signal_453 = _T_1813;
  assign rvx_signal_378 = rvx_signal_285;
  assign rvx_signal_040 = _T_1651;
  assign rvx_signal_377 = _T_1814;
  assign rvx_signal_349 = rvx_signal_087;
  assign rvx_signal_447 = _T_1656;
  assign rvx_signal_106 = _T_1815;
  assign rvx_signal_241 = rvx_signal_366;
  assign rvx_signal_078 = _T_1661;
  assign rvx_signal_134 = _T_1816;
  assign rvx_signal_365 = rvx_signal_195;
  assign rvx_signal_457 = _T_1666;
  assign rvx_signal_138 = _T_1817;
  assign rvx_signal_422 = rvx_signal_449;
  assign rvx_signal_472 = _T_1671;
  assign rvx_signal_387 = _T_1818;
  assign rvx_signal_351 = rvx_signal_363;
  assign rvx_signal_212 = _T_1676;
  assign rvx_signal_069 = _T_1819;
  assign rvx_signal_068 = rvx_signal_143;
  assign rvx_signal_473 = _T_1681;
  assign rvx_signal_160 = _T_1820;
  assign rvx_signal_118 = rvx_signal_056;
  assign rvx_signal_397 = _T_1686;
  assign rvx_signal_035 = _T_1821;
  assign rvx_signal_305 = rvx_signal_083;
  assign rvx_signal_340 = _T_1691;
  assign rvx_signal_421 = _T_1822;
  assign rvx_signal_233 = rvx_signal_314;
  assign rvx_signal_247 = _T_1696;
  assign rvx_signal_333 = _T_1823;
  assign rvx_signal_022 = rvx_signal_283;
  assign rvx_signal_274 = _T_1701;
  assign rvx_signal_020 = _T_1824;
  assign rvx_signal_086 = rvx_signal_345;
  assign rvx_signal_211 = _T_1706;
  assign rvx_signal_207 = _T_1825;
  assign rvx_signal_416 = rvx_signal_292;
  assign rvx_signal_171 = _T_1711;
  assign rvx_signal_354 = _T_1826;
  assign rvx_signal_190 = rvx_signal_136;
  assign rvx_signal_071 = _T_1716;
  assign rvx_signal_392 = _T_1827;
  assign rvx_signal_225 = rvx_signal_328;
  assign rvx_signal_094 = _T_1721;
  assign rvx_signal_176 = _T_1828;
  assign rvx_signal_469 = rvx_signal_188;
  assign rvx_signal_139 = _T_1726;
  assign rvx_signal_264 = _T_1829;
  assign rvx_signal_460 = rvx_signal_132;
  assign rvx_signal_191 = _T_1731;
  assign rvx_signal_302 = _T_1830;
  assign rvx_signal_404 = rvx_signal_406;
  assign rvx_signal_147 = _T_1736;
  assign rvx_signal_342 = _T_1831;
  assign rvx_signal_315 = rvx_signal_466;
  assign rvx_signal_105 = _T_1741;
  assign rvx_signal_467 = _T_1832;
  assign rvx_signal_003 = rvx_signal_014;
  assign rvx_signal_396 = _T_1746;
  assign rvx_signal_250 = _T_1833;
  assign rvx_signal_181 = rvx_signal_344;
  assign rvx_signal_059 = _T_1751;
  assign rvx_signal_476 = _T_1834;
  assign rvx_signal_287 = rvx_signal_208;
  assign rvx_signal_319 = _T_1756;
  assign rvx_signal_026 = _T_1835;
  assign rvx_signal_072 = rvx_signal_278;
  assign rvx_signal_260 = _T_1761;
  assign rvx_signal_478 = _T_1836;
  assign rvx_signal_276 = rvx_signal_268;
  assign rvx_signal_322 = _T_1766;
  assign rvx_signal_230 = _T_1837;
  assign rvx_signal_273 = rvx_signal_168;
  assign rvx_signal_456 = _T_1771;
  assign rvx_signal_232 = _T_1838;
  assign rvx_signal_445 = rvx_signal_196;
  assign rvx_signal_061 = _T_1776;
  assign rvx_signal_370 = _T_1839;
  assign rvx_signal_173 = rvx_signal_271;
  assign rvx_signal_286 = _T_1781;
  assign rvx_signal_339 = _T_1840;
  assign rvx_signal_189 = _T_5890;
  assign rvx_signal_161 = _T_1544;
  assign rvx_signal_017 = _T_1551;
  assign rvx_signal_164 = _T_1552;
  assign rvx_signal_427 = _T_1553;
  assign rvx_signal_005 = _T_1554;
  assign rvx_signal_275 = _T_1555;
  assign rvx_signal_182 = _T_1556;
  assign rvx_signal_185 = _T_1557;
  assign rvx_signal_110 = _T_1558;
  assign rvx_signal_372 = _T_1559;
  assign rvx_signal_290 = _T_1560;
  assign rvx_signal_407 = _T_1561;
  assign rvx_signal_126 = _T_1562;
  assign rvx_signal_374 = _T_1563;
  assign rvx_signal_318 = _T_1564;
  assign rvx_signal_279 = _T_1565;
  assign rvx_signal_303 = _T_1566;
  assign rvx_signal_038 = _T_1567;
  assign rvx_signal_077 = _T_1568;
  assign rvx_signal_384 = _T_1569;
  assign rvx_signal_446 = _T_1570;
  assign rvx_signal_443 = _T_1571;
  assign rvx_signal_150 = _T_1572;
  assign rvx_signal_383 = _T_1573;
  assign rvx_signal_048 = _T_1574;
  assign rvx_signal_249 = _T_1575;
  assign rvx_signal_064 = _T_1576;
  assign rvx_signal_470 = _T_1577;
  assign rvx_signal_258 = _T_1578;
  assign rvx_signal_034 = _T_1579;
  assign rvx_signal_018 = _T_1580;
  assign rvx_signal_155 = _T_1581;
  assign rvx_signal_144 = _T_1582;
  assign rvx_signal_431 = _T_5906;
  assign rvx_signal_120 = _T_5897;
  assign _T_1846_ready = _T_1868_ready;
  assign _T_1846_valid = _T_31_a_valid;
  assign _T_1846_bits_read = _T_1851;
  assign _T_1846_bits_index = _T_1852[23:0];
  assign _T_1846_bits_data = _T_31_a_bits_data;
  assign _T_1846_bits_mask = _T_31_a_bits_mask;
  assign _T_1846_bits_extra = _T_1853;
  assign _T_1859_ready = _T_31_d_ready;
  assign _T_1859_valid = _T_27850;
  assign _T_1859_bits_read = rvx_signal_388;
  assign _T_1859_bits_data = _T_28888;
  assign _T_1859_bits_extra = rvx_signal_263;
  assign _T_1868_ready = rvx_signal_296;
  assign _T_1868_valid = _T_1846_valid;
  assign _T_1868_bits_read = _T_1846_bits_read;
  assign _T_1868_bits_index = _T_1846_bits_index;
  assign _T_1868_bits_data = _T_1846_bits_data;
  assign _T_1868_bits_mask = _T_1846_bits_mask;
  assign _T_1868_bits_extra = _T_1846_bits_extra;
  assign rvx_signal_007 = _T_1868_valid;
  assign rvx_signal_255 = _T_1868_bits_read;
  assign rvx_signal_364 = _T_1868_bits_index;
  assign rvx_signal_129 = _T_1868_bits_data;
  assign rvx_signal_045 = _T_1868_bits_mask;
  assign rvx_signal_240 = _T_1868_bits_extra;
  assign rvx_signal_426 = _T_1859_ready;
  assign rvx_signal_043 = rvx_port_25;
  assign rvx_signal_242 = rvx_port_41;
  assign _T_3466_41 = _T_20670;
  assign _T_3573_33 = _T_23271;
  assign _T_3573_34 = _T_23311;
  assign _T_3573_35 = _T_23423;
  assign _T_3573_36 = _T_23431;
  assign _T_3573_37 = _T_23343;
  assign _T_3573_38 = _T_23391;
  assign _T_3573_39 = _T_24263;
  assign _T_3573_40 = _T_23463;
  assign _T_3573_41 = _T_25287;
  assign _T_3573_42 = _T_23239;
  assign _T_3573_43 = _T_23279;
  assign _T_3573_44 = _T_23455;
  assign _T_3573_45 = _T_23399;
  assign _T_3573_46 = _T_23303;
  assign _T_3573_47 = _T_23335;
  assign _T_3573_48 = _T_23247;
  assign _T_3573_49 = _T_23487;
  assign _T_3573_50 = _T_23367;
  assign _T_3573_51 = _T_25279;
  assign _T_3573_53 = _T_24255;
  assign _T_3573_54 = _T_24255;
  assign _T_3573_55 = _T_24255;
  assign _T_3573_56 = _T_24255;
  assign _T_3573_57 = _T_24255;
  assign _T_3573_58 = _T_24255;
  assign _T_3573_59 = _T_24255;
  assign _T_3573_60 = _T_24255;
  assign _T_3573_61 = _T_24255;
  assign _T_3573_62 = _T_24255;
  assign _T_3573_63 = _T_24255;
  assign _T_3573_64 = _T_24255;
  assign _T_3573_65 = _T_24255;
  assign _T_3573_66 = _T_24255;
  assign _T_3573_67 = _T_24255;
  assign _T_3573_68 = _T_24255;
  assign _T_3573_69 = _T_24255;
  assign _T_3573_70 = _T_24255;
  assign _T_3573_71 = _T_24255;
  assign _T_3573_72 = _T_24255;
  assign _T_3573_73 = _T_24255;
  assign _T_3573_74 = _T_24255;
  assign _T_3573_75 = _T_24255;
  assign _T_3573_76 = _T_24255;
  assign _T_3573_77 = _T_24255;
  assign _T_3573_78 = _T_24255;
  assign _T_3573_79 = _T_24255;
  assign _T_3573_80 = _T_24255;
  assign _T_3573_81 = _T_24255;
  assign _T_3573_82 = _T_24255;
  assign _T_3573_83 = _T_24255;
  assign _T_3573_84 = _T_23407;
  assign _T_3573_85 = _T_23447;
  assign _T_3573_86 = _T_23327;
  assign _T_3573_87 = _T_23287;
  assign _T_3573_88 = _T_23255;
  assign _T_3573_90 = _T_23375;
  assign _T_3573_91 = _T_23359;
  assign _T_3573_92 = _T_23479;
  assign _T_3573_93 = _T_23319;
  assign _T_3573_94 = _T_23439;
  assign _T_3573_95 = _T_23415;
  assign _T_3573_96 = _T_23295;
  assign _T_3573_97 = _T_23471;
  assign _T_3573_98 = _T_23383;
  assign _T_3573_99 = _T_23263;
  assign _T_3573_100 = _T_23351;
  assign _GEN_0 = _GEN_80;
  assign _T_27853_0 = _T_2915;
  assign _T_27853_1 = _T_3005;
  assign _T_27853_2 = _T_3059;
  assign _T_27853_3 = _T_3140;
  assign _T_27853_4 = _T_3239;
  assign _T_27853_5 = _T_2924;
  assign _T_27853_6 = _T_3014;
  assign _T_27853_7 = _T_3131;
  assign _T_27853_8 = _T_3212;
  assign _T_27853_9 = _T_3041;
  assign _T_27853_10 = _T_2933;
  assign _T_27853_11 = _T_3185;
  assign _T_27853_12 = _T_3122;
  assign _T_27853_13 = _T_3050;
  assign _T_27853_14 = _T_2960;
  assign _T_27853_15 = _T_3248;
  assign _T_27853_16 = _T_3167;
  assign _T_27853_17 = _T_3077;
  assign _T_27853_18 = _T_3158;
  assign _T_27853_19 = _T_3230;
  assign _T_27853_20 = _T_2969;
  assign _T_27853_21 = _T_3032;
  assign _T_27853_22 = _T_3104;
  assign _T_27853_23 = _T_3203;
  assign _T_27853_24 = _T_2942;
  assign _T_27853_25 = _T_2951;
  assign _T_27853_26 = _T_3194;
  assign _T_27853_27 = _T_3113;
  assign _T_27853_28 = _T_3023;
  assign _T_27853_29 = _T_2987;
  assign _T_27853_30 = _T_3221;
  assign _T_27853_31 = _T_3176;
  assign _T_27853_32 = _T_3068;
  assign _T_27853_64 = _T_2906;
  assign _T_27853_65 = _T_3149;
  assign _T_27853_128 = _T_3095;
  assign _T_27853_129 = _T_2978;
  assign _T_27853_256 = _T_3086;
  assign _T_27853_257 = _T_2996;
  assign _T_28371_1 = _T_5963;
  assign _T_28371_2 = _T_6203;
  assign _T_28371_3 = _T_7803;
  assign _T_28371_4 = _T_8243;
  assign _T_28371_5 = _T_5593;
  assign _T_28371_6 = _T_6003;
  assign _T_28371_7 = _T_7763;
  assign _T_28371_8 = _T_8123;
  assign _T_28371_9 = _T_6123;
  assign _T_28371_10 = _T_5633;
  assign _T_28371_11 = _T_8003;
  assign _T_28371_12 = _T_7723;
  assign _T_28371_13 = _T_6163;
  assign _T_28371_14 = _T_5753;
  assign _T_28371_15 = _T_8283;
  assign _T_28371_16 = _T_7923;
  assign _T_28371_17 = _T_6283;
  assign _T_28371_18 = _T_7883;
  assign _T_28371_19 = _T_8203;
  assign _T_28371_20 = _T_5793;
  assign _T_28371_21 = _T_6083;
  assign _T_28371_22 = _T_7643;
  assign _T_28371_23 = _T_8083;
  assign _T_28371_24 = _T_5673;
  assign _T_28371_25 = _T_5713;
  assign _T_28371_26 = _T_8043;
  assign _T_28371_27 = _T_7683;
  assign _T_28371_28 = _T_6043;
  assign _T_28371_29 = _T_5873;
  assign _T_28371_30 = _T_8163;
  assign _T_28371_31 = _T_7963;
  assign _T_28371_32 = _T_6243;
  assign _T_28371_64 = _T_5514;
  assign _T_28371_65 = {{31'd0}, rvx_signal_229};
  assign _T_28371_128 = _T_7604;
  assign _T_28371_129 = {{31'd0}, rvx_signal_408};
  assign _T_28371_256 = _T_6323;
  assign _T_28371_257 = _T_5923;
  assign _GEN_5 = _GEN_2693;
  assign _GEN_6 = _GEN_3204;
  assign _T_28893_size = _T_28890;
  assign _T_28893_source = _T_28889;

always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_243 <= 0;
  end
  else
    rvx_signal_243 <= _GEN_81[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_057 <= 0;
  end
  else
    rvx_signal_057 <= _GEN_87[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_311 <= 0;
  end
  else
    rvx_signal_311 <= _GEN_127[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_089 <= 0;
  end
  else
    rvx_signal_089 <= _GEN_137[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_117 <= 0;
  end
  else
    rvx_signal_117 <= _GEN_41[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_116 <= 0;
  end
  else
    rvx_signal_116 <= _GEN_82[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_415 <= 0;
  end
  else
    rvx_signal_415 <= _GEN_126[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_289 <= 0;
  end
  else
    rvx_signal_289 <= _GEN_134[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_002 <= 0;
  end
  else
    rvx_signal_002 <= _GEN_85[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_395 <= 0;
  end
  else
    rvx_signal_395 <= _GEN_42[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_140 <= 0;
  end
  else
    rvx_signal_140 <= _GEN_131[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_023 <= 0;
  end
  else
    rvx_signal_023 <= _GEN_125[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_145 <= 0;
  end
  else
    rvx_signal_145 <= _GEN_86[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_025 <= 0;
  end
  else
    rvx_signal_025 <= _GEN_45[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_418 <= 0;
  end
  else
    rvx_signal_418 <= _GEN_138[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_008 <= 0;
  end
  else
    rvx_signal_008 <= _GEN_129[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_245 <= 0;
  end
  else
    rvx_signal_245 <= _GEN_89[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_114 <= 0;
  end
  else
    rvx_signal_114 <= _GEN_128[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_172 <= 0;
  end
  else
    rvx_signal_172 <= _GEN_136[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_266 <= 0;
  end
  else
    rvx_signal_266 <= _GEN_46[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_444 <= 0;
  end
  else
    rvx_signal_444 <= _GEN_84[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_088 <= 0;
  end
  else
    rvx_signal_088 <= _GEN_123[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_234 <= 0;
  end
  else
    rvx_signal_234 <= _GEN_133[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_097 <= 0;
  end
  else
    rvx_signal_097 <= _GEN_43[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_267 <= 0;
  end
  else
    rvx_signal_267 <= _GEN_44[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_248 <= 0;
  end
  else
    rvx_signal_248 <= _GEN_132[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_400 <= 0;
  end
  else
    rvx_signal_400 <= _GEN_124[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_430 <= 0;
  end
  else
    rvx_signal_430 <= _GEN_83[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_359 <= 0;
  end
  else
    rvx_signal_359 <= _GEN_48[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_332 <= 0;
  end
  else
    rvx_signal_332 <= _GEN_135[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_300 <= 0;
  end
  else
    rvx_signal_300 <= _GEN_130[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_032 <= 0;
  end
  else
    rvx_signal_032 <= _GEN_88[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_435 <= 0;
  end
  else
    rvx_signal_435 <= _GEN_90[2:0];
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_065 <= 1'h0;
  end else begin
    if (_T_1627) begin
      rvx_signal_065 <= _T_1629;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_437 <= 1'h0;
  end else begin
    if (_T_1632) begin
      rvx_signal_437 <= _T_1634;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_382 <= 1'h0;
  end else begin
    if (_T_1637) begin
      rvx_signal_382 <= _T_1639;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_316 <= 1'h0;
  end else begin
    if (_T_1642) begin
      rvx_signal_316 <= _T_1644;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_165 <= 1'h0;
  end else begin
    if (_T_1647) begin
      rvx_signal_165 <= _T_1649;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_004 <= 1'h0;
  end else begin
    if (_T_1652) begin
      rvx_signal_004 <= _T_1654;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_272 <= 1'h0;
  end else begin
    if (_T_1657) begin
      rvx_signal_272 <= _T_1659;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_409 <= 1'h0;
  end else begin
    if (_T_1662) begin
      rvx_signal_409 <= _T_1664;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_202 <= 1'h0;
  end else begin
    if (_T_1667) begin
      rvx_signal_202 <= _T_1669;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_454 <= 1'h0;
  end else begin
    if (_T_1672) begin
      rvx_signal_454 <= _T_1674;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_092 <= 1'h0;
  end else begin
    if (_T_1677) begin
      rvx_signal_092 <= _T_1679;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_298 <= 1'h0;
  end else begin
    if (_T_1682) begin
      rvx_signal_298 <= _T_1684;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_096 <= 1'h0;
  end else begin
    if (_T_1687) begin
      rvx_signal_096 <= _T_1689;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_167 <= 1'h0;
  end else begin
    if (_T_1692) begin
      rvx_signal_167 <= _T_1694;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_294 <= 1'h0;
  end else begin
    if (_T_1697) begin
      rvx_signal_294 <= _T_1699;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_371 <= 1'h0;
  end else begin
    if (_T_1702) begin
      rvx_signal_371 <= _T_1704;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_103 <= 1'h0;
  end else begin
    if (_T_1707) begin
      rvx_signal_103 <= _T_1709;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_019 <= 1'h0;
  end else begin
    if (_T_1712) begin
      rvx_signal_019 <= _T_1714;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_080 <= 1'h0;
  end else begin
    if (_T_1717) begin
      rvx_signal_080 <= _T_1719;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_239 <= 1'h0;
  end else begin
    if (_T_1722) begin
      rvx_signal_239 <= _T_1724;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_124 <= 1'h0;
  end else begin
    if (_T_1727) begin
      rvx_signal_124 <= _T_1729;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_222 <= 1'h0;
  end else begin
    if (_T_1732) begin
      rvx_signal_222 <= _T_1734;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_306 <= 1'h0;
  end else begin
    if (_T_1737) begin
      rvx_signal_306 <= _T_1739;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_238 <= 1'h0;
  end else begin
    if (_T_1742) begin
      rvx_signal_238 <= _T_1744;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_011 <= 1'h0;
  end else begin
    if (_T_1747) begin
      rvx_signal_011 <= _T_1749;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_029 <= 1'h0;
  end else begin
    if (_T_1752) begin
      rvx_signal_029 <= _T_1754;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_166 <= 1'h0;
  end else begin
    if (_T_1757) begin
      rvx_signal_166 <= _T_1759;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_228 <= 1'h0;
  end else begin
    if (_T_1762) begin
      rvx_signal_228 <= _T_1764;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_183 <= 1'h0;
  end else begin
    if (_T_1767) begin
      rvx_signal_183 <= _T_1769;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_253 <= 1'h0;
  end else begin
    if (_T_1772) begin
      rvx_signal_253 <= _T_1774;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_033 <= 1'h0;
  end else begin
    if (_T_1777) begin
      rvx_signal_033 <= _T_1779;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_229 <= 1'h0;
  end else begin
    if (_T_1782) begin
      rvx_signal_229 <= _T_1784;
    end
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_099 <= 0;
  end
  else if (_T_6384) begin
    rvx_signal_099 <= _T_4295;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_369 <= 0;
  end
  else if (_T_6424) begin
    rvx_signal_369 <= _T_4335;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_221 <= 0;
  end
  else if (_T_6464) begin
    rvx_signal_221 <= _T_4375;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_224 <= 0;
  end
  else if (_T_6504) begin
    rvx_signal_224 <= _T_4415;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_066 <= 0;
  end
  else if (_T_6544) begin
    rvx_signal_066 <= _T_4455;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_111 <= 0;
  end
  else if (_T_6584) begin
    rvx_signal_111 <= _T_4495;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_179 <= 0;
  end
  else if (_T_6624) begin
    rvx_signal_179 <= _T_4535;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_050 <= 0;
  end
  else if (_T_6664) begin
    rvx_signal_050 <= _T_4575;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_215 <= 0;
  end
  else if (_T_6704) begin
    rvx_signal_215 <= _T_4615;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_386 <= 0;
  end
  else if (_T_6744) begin
    rvx_signal_386 <= _T_4655;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_450 <= 0;
  end
  else if (_T_6784) begin
    rvx_signal_450 <= _T_4695;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_399 <= 0;
  end
  else if (_T_6824) begin
    rvx_signal_399 <= _T_4735;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_067 <= 0;
  end
  else if (_T_6864) begin
    rvx_signal_067 <= _T_4775;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_350 <= 0;
  end
  else if (_T_6904) begin
    rvx_signal_350 <= _T_4815;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_265 <= 0;
  end
  else if (_T_6944) begin
    rvx_signal_265 <= _T_4855;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_304 <= 0;
  end
  else if (_T_6984) begin
    rvx_signal_304 <= _T_4895;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_058 <= 0;
  end
  else if (_T_7024) begin
    rvx_signal_058 <= _T_4935;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_433 <= 0;
  end
  else if (_T_7064) begin
    rvx_signal_433 <= _T_4975;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_465 <= 0;
  end
  else if (_T_7104) begin
    rvx_signal_465 <= _T_5015;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_197 <= 0;
  end
  else if (_T_7144) begin
    rvx_signal_197 <= _T_5055;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_358 <= 0;
  end
  else if (_T_7184) begin
    rvx_signal_358 <= _T_5095;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_436 <= 0;
  end
  else if (_T_7224) begin
    rvx_signal_436 <= _T_5135;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_001 <= 0;
  end
  else if (_T_7264) begin
    rvx_signal_001 <= _T_5175;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_131 <= 0;
  end
  else if (_T_7304) begin
    rvx_signal_131 <= _T_5215;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_410 <= 0;
  end
  else if (_T_7344) begin
    rvx_signal_410 <= _T_5255;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_137 <= 0;
  end
  else if (_T_7384) begin
    rvx_signal_137 <= _T_5295;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_178 <= 0;
  end
  else if (_T_7424) begin
    rvx_signal_178 <= _T_5335;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_052 <= 0;
  end
  else if (_T_7464) begin
    rvx_signal_052 <= _T_5375;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_423 <= 0;
  end
  else if (_T_7504) begin
    rvx_signal_423 <= _T_5415;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_462 <= 0;
  end
  else if (_T_7544) begin
    rvx_signal_462 <= _T_5455;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_475 <= 0;
  end
  else if (_T_7584) begin
    rvx_signal_475 <= _T_5495;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_408 <= 0;
  end
  else if (_T_5814) begin
    rvx_signal_408 <= _T_4255;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    rvx_signal_153 <= 0;
  end
  else if (_T_1511) begin
    rvx_signal_153 <= {{1'd0}, _T_1509};
  end else begin
    rvx_signal_153 <= 6'h20;
  end
end
always @(posedge rvx_port_25, posedge rvx_port_41) begin
  if (rvx_port_41) begin
    _T_1517 <= 0;
  end
  else if (_T_1511) begin
    if (_T_1505) begin
      if (_T_1409) begin
        if (_T_1361) begin
          if (_T_1337) begin
            if (_T_1325) begin
              _T_1517 <= 4'h8;
            end else begin
              _T_1517 <= _T_1260;
            end
          end else begin
            if (_T_1332) begin
              _T_1517 <= _T_1262;
            end else begin
              _T_1517 <= _T_1264;
            end
          end
        end else begin
          if (_T_1356) begin
            if (_T_1344) begin
              _T_1517 <= _T_1266;
            end else begin
              _T_1517 <= _T_1268;
            end
          end else begin
            if (_T_1351) begin
              _T_1517 <= _T_1270;
            end else begin
              _T_1517 <= _T_1272;
            end
          end
        end
      end else begin
        if (_T_1404) begin
          if (_T_1380) begin
            if (_T_1368) begin
              _T_1517 <= _T_1274;
            end else begin
              _T_1517 <= _T_1276;
            end
          end else begin
            if (_T_1375) begin
              _T_1517 <= _T_1278;
            end else begin
              _T_1517 <= _T_1280;
            end
          end
        end else begin
          if (_T_1399) begin
            if (_T_1387) begin
              _T_1517 <= _T_1282;
            end else begin
              _T_1517 <= _T_1284;
            end
          end else begin
            if (_T_1394) begin
              _T_1517 <= _T_1286;
            end else begin
              _T_1517 <= _T_1288;
            end
          end
        end
      end
    end else begin
      if (_T_1500) begin
        if (_T_1452) begin
          if (_T_1428) begin
            if (_T_1416) begin
              _T_1517 <= _T_1290;
            end else begin
              _T_1517 <= _T_1292;
            end
          end else begin
            if (_T_1423) begin
              _T_1517 <= _T_1294;
            end else begin
              _T_1517 <= _T_1296;
            end
          end
        end else begin
          if (_T_1447) begin
            if (_T_1435) begin
              _T_1517 <= _T_1298;
            end else begin
              _T_1517 <= _T_1300;
            end
          end else begin
            if (_T_1442) begin
              _T_1517 <= _T_1302;
            end else begin
              _T_1517 <= _T_1304;
            end
          end
        end
      end else begin
        if (_T_1495) begin
          if (_T_1471) begin
            if (_T_1459) begin
              _T_1517 <= _T_1306;
            end else begin
              _T_1517 <= _T_1308;
            end
          end else begin
            if (_T_1466) begin
              _T_1517 <= _T_1310;
            end else begin
              _T_1517 <= _T_1312;
            end
          end
        end else begin
          if (_T_1490) begin
            if (_T_1478) begin
              _T_1517 <= _T_1314;
            end else begin
              _T_1517 <= _T_1316;
            end
          end else begin
            if (_T_1485) begin
              _T_1517 <= _T_1318;
            end else begin
              _T_1517 <= _T_1320;
            end
          end
        end
      end
    end
  end else begin
    _T_1517 <= _T_1322;
  end
end
endmodule
