
/*****************************************************************************
 *
 * Copyright Embedded DSP Development Group 2006-2009, All rights reserved.
 * Electronics and Telecommunications Research Institute (ETRI)
 *
 * THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE 
 * WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS 
 * TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE REPRODUCED, 
 * COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL SYSTEM OR 
 * TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE, IN ANY FORM, 
 * BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE COMPLETE PRIOR WRITTEN 
 * PERMISSION OF ETRI.
 *
 *****************************************************************************
 *
 * UART macro definitions
 *
 *****************************************************************************/


//--------------------------------------------------------------------
// UART Internal SFR definitions
//--------------------------------------------------------------------
//(Note) The following defintions are replaced statically.
//`define __ERVP_UART_DEFINES_H__
//`define UART_DATA_WIDTH 8
//`define UART_HAS_BAUDRATE_OUTPUT

`include "ervp_misc_util.vh"
`include "platform_info.vh"

`define UART_ADDR_DIFF 8
`define BW_UART_REG_INDEX (4+`PLOG2(`UART_ADDR_DIFF))

// Register addresses
`define UART_REG_RB		(0*`UART_ADDR_DIFF)	// receiver buffer
`define UART_REG_TR  	(0*`UART_ADDR_DIFF) // transmitter
`define UART_REG_IE		(1*`UART_ADDR_DIFF)	// Interrupt enable
`define UART_REG_II  	(2*`UART_ADDR_DIFF)	// Interrupt identification
`define UART_REG_FC  	(2*`UART_ADDR_DIFF) // FIFO control
`define UART_REG_LC		(3*`UART_ADDR_DIFF) // Line Control
`define UART_REG_MC		(4*`UART_ADDR_DIFF) // Modem control
`define UART_REG_LS  	(5*`UART_ADDR_DIFF) // Line status
`define UART_REG_MS  	(6*`UART_ADDR_DIFF) // Modem status
`define UART_REG_SR  	(7*`UART_ADDR_DIFF) // Scratch register
`define UART_REG_EN  	(8*`UART_ADDR_DIFF) // UART Enable
`define UART_REG_TC  	(9*`UART_ADDR_DIFF) // tranmitter count

`define UART_REG_DL1	(4'd0)	// Divisor latch bytes (1-2)
`define UART_REG_DL2	(4'd1)

// Interrupt Enable register bits
`define UART_IE_RDA		0	// Received Data available interrupt
`define UART_IE_THRE	1	// Transmitter Holding Register empty interrupt
`define UART_IE_RLS		2	// Receiver Line Status Interrupt
`define UART_IE_MS		3	// Modem Status Interrupt

// Interrupt Identification register bits
`define UART_II_IP		0	// Interrupt pending when 0
`define UART_II_II		3:1	// Interrupt identification

// Interrupt identification values for bits 3:1
`define UART_II_RLS		3'b011	// Receiver Line Status
`define UART_II_RDA		3'b010	// Receiver Data available
`define UART_II_TI		3'b110	// Timeout Indication
`define UART_II_THRE	3'b001	// Transmitter Holding Register empty
`define UART_II_MS		3'b000	// Modem Status

// FIFO Control Register bits
`define UART_FC_TL		1:0	// Trigger level

// FIFO trigger level values
`define UART_FC_1		2'b00
`define UART_FC_4		2'b01
`define UART_FC_8		2'b10
`define UART_FC_14		2'b11

// Line Control register bits
`define UART_LC_BITS	1:0	// bits in character
`define UART_LC_SB		2	// stop bits
`define UART_LC_PE		3	// parity enable
`define UART_LC_EP		4	// even parity
`define UART_LC_SP		5	// stick parity
`define UART_LC_BC		6	// Break control
`define UART_LC_DL		7	// Divisor Latch access bit

// Modem Control register bits
`define UART_MC_DTR		0
`define UART_MC_RTS		1
`define UART_MC_OUT1	2
`define UART_MC_OUT2	3
`define UART_MC_LB	4	// Loopback mode

// Line Status Register bits
`define UART_LS_DR		0	// Data ready
`define UART_LS_OE		1	// Overrun Error
`define UART_LS_PE		2	// Parity Error
`define UART_LS_FE		3	// Framing Error
`define UART_LS_BI		4	// Break interrupt
`define UART_LS_TFE		5	// Transmit FIFO is empty
`define UART_LS_TE		6	// Transmitter Empty indicator
`define UART_LS_EI		7	// Error indicator

// Modem Status Register bits
`define UART_MS_DCTS	0	// Delta signals
`define UART_MS_DDSR	1
`define UART_MS_TERI	2
`define UART_MS_DDCD	3
`define UART_MS_CCTS	4	// Complement signals
`define UART_MS_CDSR	5
`define UART_MS_CRI		6
`define UART_MS_CDCD	7

// FIFO parameter defines

`define UART_FIFO_WIDTH		8

`ifndef UART_FIFO_DEPTH
`define UART_FIFO_DEPTH 128
`endif

// receiver fifo has width 11 because it has break, parity and framing error bits
`define UART_FIFO_REC_WIDTH  11

