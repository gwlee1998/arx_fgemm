// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_227
`define RVX_GDEF_227

`define RVX_GDEF_281 8
`define RVX_GDEF_124 8
`define RVX_GDEF_285 3
`define RVX_GDEF_195 1

`define RVX_GDEF_396 (32'h 0)
`define RVX_GDEF_303 (32'h 8)
`define RVX_GDEF_068 (32'h 10)
`define RVX_GDEF_245 (32'h 18)
`define RVX_GDEF_223 (32'h 20)
`define RVX_GDEF_314 (32'h 28)
`define RVX_GDEF_292 (32'h 30)
`define RVX_GDEF_009 (32'h 38)
`define RVX_GDEF_013 (32'h 40)
`define RVX_GDEF_394 (32'h 48)
`define RVX_GDEF_432 (32'h 50)
`define RVX_GDEF_324 (32'h 58)
`define RVX_GDEF_265 (32'h 60)
`define RVX_GDEF_371 (32'h 68)
`define RVX_GDEF_225 (32'h 70)
`define RVX_GDEF_169 (32'h 78)
`define RVX_GDEF_005 (32'h 80)
`define RVX_GDEF_251 (32'h 88)
`define RVX_GDEF_435 (32'h 90)
`define RVX_GDEF_180 (32'h 98)
`define RVX_GDEF_115 (32'h a0)
`define RVX_GDEF_163 (32'h a8)
`define RVX_GDEF_295 (32'h b0)
`define RVX_GDEF_244 (32'h b8)
`define RVX_GDEF_107 (32'h c0)

`define RVX_GDEF_316 (`RVX_GDEF_396)
`define RVX_GDEF_166 (`RVX_GDEF_303)
`define RVX_GDEF_192 (`RVX_GDEF_068)
`define RVX_GDEF_079 (`RVX_GDEF_245)
`define RVX_GDEF_047 (`RVX_GDEF_223)
`define RVX_GDEF_317 (`RVX_GDEF_314)
`define RVX_GDEF_172 (`RVX_GDEF_292)
`define RVX_GDEF_145 (`RVX_GDEF_009)
`define RVX_GDEF_367 (`RVX_GDEF_013)
`define RVX_GDEF_349 (`RVX_GDEF_394)
`define RVX_GDEF_055 (`RVX_GDEF_432)
`define RVX_GDEF_089 (`RVX_GDEF_324)
`define RVX_GDEF_038 (`RVX_GDEF_265)
`define RVX_GDEF_372 (`RVX_GDEF_371)
`define RVX_GDEF_420 (`RVX_GDEF_225)
`define RVX_GDEF_388 (`RVX_GDEF_169)
`define RVX_GDEF_397 (`RVX_GDEF_005)
`define RVX_GDEF_074 (`RVX_GDEF_251)
`define RVX_GDEF_364 (`RVX_GDEF_435)
`define RVX_GDEF_203 (`RVX_GDEF_180)
`define RVX_GDEF_284 (`RVX_GDEF_115)
`define RVX_GDEF_264 (`RVX_GDEF_163)
`define RVX_GDEF_333 (`RVX_GDEF_295)
`define RVX_GDEF_143 (`RVX_GDEF_244)
`define RVX_GDEF_114 (`RVX_GDEF_107)

`define RVX_GDEF_036 8
`define RVX_GDEF_049 0

`define RVX_GDEF_290 32
`define RVX_GDEF_377 0

`define RVX_GDEF_185 32
`define RVX_GDEF_031 0

`define RVX_GDEF_088 32
`define RVX_GDEF_408 0

`endif