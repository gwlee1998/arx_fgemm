`ifndef __DCA_MATRIX_QGEMM_DEFINES_H__
`define __DCA_MATRIX_QGEMM_DEFINES_H__

`define BW_DCA_MATRIX_QDQ_INST 512
`define DCA_MATRIX_QDQ_INST_DEFAULT_VALUE 0

`define BW_DCA_MATRIX_QDQ_LOG 32
`define DCA_MATRIX_QDQ_LOG_DEFAULT_VALUE 0

`define BW_DCA_MATRIX_QDQ_STATUS 32
`define DCA_MATRIX_QDQ_STATUS_DEFAULT_VALUE 0

`define DCA_MATRIX_QDQ_NUM_COL 16
`define DCA_MATRIX_QDQ_NUM_ROW 16
`define QUANT_PRECCISION_NUM_BIT 8

`define QUANT_USING_EXP_AND_MANTISSA 1
// `define QUANT_USING_ONLY_EXP
`define USE_OPT_QUANT 1

`endif

