// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_158
`define RVX_GDEF_158

`define RVX_GDEF_016 6
`define RVX_GDEF_390 8
`define RVX_GDEF_004 3
`define RVX_GDEF_370 1

`define RVX_GDEF_224 (32'h 0)
`define RVX_GDEF_287 (32'h 8)
`define RVX_GDEF_386 (32'h 10)
`define RVX_GDEF_311 (32'h 18)
`define RVX_GDEF_325 (32'h 20)
`define RVX_GDEF_354 (32'h 28)

`define RVX_GDEF_312 (`RVX_GDEF_224)
`define RVX_GDEF_252 (`RVX_GDEF_287)
`define RVX_GDEF_299 (`RVX_GDEF_386)
`define RVX_GDEF_253 (`RVX_GDEF_311)
`define RVX_GDEF_437 (`RVX_GDEF_325)
`define RVX_GDEF_286 (`RVX_GDEF_354)

`define RVX_GDEF_018 8
`define RVX_GDEF_102 0
`define RVX_GDEF_300 1
`define RVX_GDEF_043 2
`define RVX_GDEF_352 4
`define RVX_GDEF_326 8
`define RVX_GDEF_092 16
`define RVX_GDEF_012 32
`define RVX_GDEF_148 64
`define RVX_GDEF_320 128
`define RVX_GDEF_379 0
`define RVX_GDEF_177 1
`define RVX_GDEF_419 2
`define RVX_GDEF_023 3
`define RVX_GDEF_046 4
`define RVX_GDEF_008 5
`define RVX_GDEF_168 6
`define RVX_GDEF_240 7
`define RVX_GDEF_250 0

`define RVX_GDEF_260 5
`define RVX_GDEF_206 0
`define RVX_GDEF_099 1
`define RVX_GDEF_215 2
`define RVX_GDEF_234 4
`define RVX_GDEF_035 8
`define RVX_GDEF_188 16
`define RVX_GDEF_366 0
`define RVX_GDEF_288 1
`define RVX_GDEF_330 2
`define RVX_GDEF_041 3
`define RVX_GDEF_258 4
`define RVX_GDEF_263 0

`define RVX_GDEF_318 8
`define RVX_GDEF_056 0

`define RVX_GDEF_161 32
`define RVX_GDEF_211 0

`define RVX_GDEF_003 32
`define RVX_GDEF_123 0

`define RVX_GDEF_332 7
`define RVX_GDEF_369 0

`endif