// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************

localparam MMIOX1_FIFO_PARA_0_AFTER = MMIOX1_FIFO_PARA;

localparam MMIOX1_FIFO_PARA_1_ANDSOON = MMIOX1_FIFO_PARA_0_AFTER;
localparam MMIOX1_FIFO_PARA_1_AFTER = MMIOX1_FIFO_PARA_1_ANDSOON >> MMIOX1_FIFO_PARA_1_BIT;
localparam _LOG_FIFO_DEPTH_TEMP = MMIOX1_FIFO_PARA_1_ANDSOON % (2**MMIOX1_FIFO_PARA_1_BIT);
localparam INCLUDE_LOG_FIFO = (_LOG_FIFO_DEPTH_TEMP!=0);
localparam LOG_FIFO_DEPTH = `MAX(2, _LOG_FIFO_DEPTH_TEMP);
localparam LOG_FIFO_DEPTH_DEFAULT = 4;

localparam MMIOX1_FIFO_PARA_2_ANDSOON = MMIOX1_FIFO_PARA_1_AFTER;
localparam MMIOX1_FIFO_PARA_2_AFTER = MMIOX1_FIFO_PARA_2_ANDSOON >> MMIOX1_FIFO_PARA_2_BIT;
localparam _INST_FIFO_DEPTH_TEMP = MMIOX1_FIFO_PARA_2_ANDSOON % (2**MMIOX1_FIFO_PARA_2_BIT);
localparam INCLUDE_INST_FIFO = (_INST_FIFO_DEPTH_TEMP!=0);
localparam INST_FIFO_DEPTH = `MAX(2, _INST_FIFO_DEPTH_TEMP);
localparam INST_FIFO_DEPTH_DEFAULT = 4;

localparam MMIOX1_FIFO_PARA_3_ANDSOON = MMIOX1_FIFO_PARA_2_AFTER;
localparam MMIOX1_FIFO_PARA_3_AFTER = MMIOX1_FIFO_PARA_3_ANDSOON >> MMIOX1_FIFO_PARA_3_BIT;
localparam _INPUT_FIFO_DEPTH_TEMP = MMIOX1_FIFO_PARA_3_ANDSOON % (2**MMIOX1_FIFO_PARA_3_BIT);
localparam INCLUDE_INPUT_FIFO = (_INPUT_FIFO_DEPTH_TEMP!=0);
localparam INPUT_FIFO_DEPTH = `MAX(2, _INPUT_FIFO_DEPTH_TEMP);
localparam INPUT_FIFO_DEPTH_DEFAULT = 4;

localparam MMIOX1_FIFO_PARA_4_ANDSOON = MMIOX1_FIFO_PARA_3_AFTER;
localparam MMIOX1_FIFO_PARA_4_AFTER = MMIOX1_FIFO_PARA_4_ANDSOON >> MMIOX1_FIFO_PARA_4_BIT;
localparam _OUTPUT_FIFO_DEPTH_TEMP = MMIOX1_FIFO_PARA_4_ANDSOON % (2**MMIOX1_FIFO_PARA_4_BIT);
localparam INCLUDE_OUTPUT_FIFO = (_OUTPUT_FIFO_DEPTH_TEMP!=0);
localparam OUTPUT_FIFO_DEPTH = `MAX(2, _OUTPUT_FIFO_DEPTH_TEMP);
localparam OUTPUT_FIFO_DEPTH_DEFAULT = 4;
