`ifndef __ERVP_TRIGGER_COND_MEMORYMAP_OFFSET_H__
`define __ERVP_TRIGGER_COND_MEMORYMAP_OFFSET_H__



// reg ervp_trigger_cond
`define BW_ERVP_TRIGGER_COND 5
`define ERVP_TRIGGER_COND_DEFAULT_VALUE 0
`define ERVP_TRIGGER_COND_HIGH 1
`define ERVP_TRIGGER_COND_LOW 2
`define ERVP_TRIGGER_COND_RISE 4
`define ERVP_TRIGGER_COND_FALL 8
`define ERVP_TRIGGER_COND_EQ 16
`define ERVP_TRIGGER_COND_INDEX_HIGH 0
`define ERVP_TRIGGER_COND_INDEX_LOW 1
`define ERVP_TRIGGER_COND_INDEX_RISE 2
`define ERVP_TRIGGER_COND_INDEX_FALL 3
`define ERVP_TRIGGER_COND_INDEX_EQ 4
`define ERVP_TRIGGER_COND_NONE 0

`endif