// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL 
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE, 
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE 
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2019-03
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************

`ifndef __MUNOC_NETWORK_INCLUDE_H__
`define __MUNOC_NETWORK_INCLUDE_H__

`include "munoc_include_04.vh"
`include "munoc_extended_config.vh"
`include "munoc_network_type.vh"
`include "munoc_network_link.vh"
`include "munoc_arbitration_type.vh"
`include "munoc_tid_control_type.vh"
`include "munoc_include_10.vh"
`include "munoc_control.vh"
`include "ervp_axi_define.vh"
`include "ervp_ahb_define.vh"

`include "munoc_node_id.vh"
`include "munoc_router_id.vh"
`include "munoc_process_id.vh"

`endif
