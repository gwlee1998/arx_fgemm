// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_436
`define RVX_GDEF_436

`define RVX_GDEF_389 15
`define RVX_GDEF_319 8
`define RVX_GDEF_184 3
`define RVX_GDEF_327 6
`define RVX_GDEF_310 3
`define RVX_GDEF_159 0
`define RVX_GDEF_382 (32'h 0)
`define RVX_GDEF_410 1
`define RVX_GDEF_343 (32'h 1000)
`define RVX_GDEF_063 2
`define RVX_GDEF_413 (32'h 2000)
`define RVX_GDEF_131 3
`define RVX_GDEF_231 (32'h 3000)
`define RVX_GDEF_026 4
`define RVX_GDEF_085 (32'h 4000)
`define RVX_GDEF_296 5
`define RVX_GDEF_351 (32'h 5000)

`define RVX_GDEF_073 8
`define RVX_GDEF_280 3

`define RVX_GDEF_173 5
`define RVX_GDEF_315 3
`define RVX_GDEF_368 (32'h 0)
`define RVX_GDEF_363 (32'h 8)
`define RVX_GDEF_307 (32'h 10)

`define RVX_GDEF_170 (`RVX_GDEF_343+`RVX_GDEF_368)
`define RVX_GDEF_236 (`RVX_GDEF_343+`RVX_GDEF_363)
`define RVX_GDEF_407 (`RVX_GDEF_343+`RVX_GDEF_307)

`define RVX_GDEF_338 12
`define RVX_GDEF_270 3

`define RVX_GDEF_269 10
`define RVX_GDEF_405 3

`define RVX_GDEF_361 10
`define RVX_GDEF_164 3

`define RVX_GDEF_248 8
`define RVX_GDEF_104 3

`define RVX_GDEF_309 8
`define RVX_GDEF_339 0

`define RVX_GDEF_030 8
`define RVX_GDEF_404 0

`define RVX_GDEF_120 1
`define RVX_GDEF_066 0

`endif