// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_336
`define RVX_GDEF_336

`define RVX_GDEF_101 5
`define RVX_GDEF_083 8
`define RVX_GDEF_132 3
`define RVX_GDEF_308 1

`define RVX_GDEF_077 (32'h 0)
`define RVX_GDEF_080 (32'h 8)
`define RVX_GDEF_078 (32'h 10)

`define RVX_GDEF_028 (`RVX_GDEF_077)
`define RVX_GDEF_294 (`RVX_GDEF_080)
`define RVX_GDEF_126 (`RVX_GDEF_078)

`define RVX_GDEF_238 32
`define RVX_GDEF_301 0

`define RVX_GDEF_346 32
`define RVX_GDEF_154 0

`define RVX_GDEF_067 2
`define RVX_GDEF_204 0

`define RVX_GDEF_133 5
`define RVX_GDEF_149 0
`define RVX_GDEF_232 1
`define RVX_GDEF_212 2
`define RVX_GDEF_200 4
`define RVX_GDEF_040 8
`define RVX_GDEF_358 16
`define RVX_GDEF_072 0
`define RVX_GDEF_282 1
`define RVX_GDEF_403 2
`define RVX_GDEF_378 3
`define RVX_GDEF_157 4
`define RVX_GDEF_293 0

`define RVX_GDEF_360 2
`define RVX_GDEF_086 0
`define RVX_GDEF_019 0
`define RVX_GDEF_267 1
`define RVX_GDEF_002 2
`define RVX_GDEF_249 3
`define RVX_GDEF_289 0
`define RVX_GDEF_218 1

`define RVX_GDEF_001 3
`define RVX_GDEF_230 0
`define RVX_GDEF_247 0
`define RVX_GDEF_112 1
`define RVX_GDEF_135 2
`define RVX_GDEF_141 3
`define RVX_GDEF_305 4
`define RVX_GDEF_090 5
`define RVX_GDEF_011 0
`define RVX_GDEF_323 1
`define RVX_GDEF_060 2

`endif