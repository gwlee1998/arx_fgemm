`default_nettype wire
`include "timescale.vh"
module FPUDecoder(
  input  [31:0] io_inst,
  output        io_sigs_wen,
  output        io_sigs_ren1,
  output        io_sigs_ren2,
  output        io_sigs_ren3,
  output        io_sigs_swap12,
  output        io_sigs_swap23,
  output [1:0]  io_sigs_typeTagOut,
  output        io_sigs_fromint,
  output        io_sigs_toint,
  output        io_sigs_fastpipe,
  output        io_sigs_fma,
  output        io_sigs_div,
  output        io_sigs_sqrt,
  output        io_sigs_wflags
);
  wire [31:0] decoder_decoded_invInputs = ~io_inst;
  wire  decoder_decoded_andMatrixInput_0 = io_inst[0];
  wire  decoder_decoded_andMatrixInput_1 = io_inst[1];
  wire  decoder_decoded_andMatrixInput_2 = decoder_decoded_invInputs[4];
  wire  decoder_decoded_andMatrixInput_3 = decoder_decoded_invInputs[5];
  wire  decoder_decoded_andMatrixInput_4 = io_inst[6];
  wire [4:0] _decoder_decoded_T = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2,decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4};
  wire  _decoder_decoded_T_1 = &_decoder_decoded_T;
  wire  decoder_decoded_andMatrixInput_2_1 = decoder_decoded_invInputs[2];
  wire  decoder_decoded_andMatrixInput_3_1 = decoder_decoded_invInputs[3];
  wire  decoder_decoded_andMatrixInput_4_1 = io_inst[4];
  wire  decoder_decoded_andMatrixInput_7 = decoder_decoded_invInputs[25];
  wire  decoder_decoded_andMatrixInput_8 = decoder_decoded_invInputs[26];
  wire  decoder_decoded_andMatrixInput_9 = decoder_decoded_invInputs[29];
  wire  decoder_decoded_andMatrixInput_10 = decoder_decoded_invInputs[30];
  wire  decoder_decoded_andMatrixInput_11 = decoder_decoded_invInputs[31];
  wire [5:0] decoder_decoded_lo_1 = {decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9,decoder_decoded_andMatrixInput_10,
    decoder_decoded_andMatrixInput_11};
  wire [11:0] _decoder_decoded_T_2 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_lo_1};
  wire  _decoder_decoded_T_3 = &_decoder_decoded_T_2;
  wire  decoder_decoded_andMatrixInput_9_1 = decoder_decoded_invInputs[27];
  wire [5:0] decoder_decoded_lo_2 = {decoder_decoded_andMatrixInput_7,decoder_decoded_andMatrixInput_8,
    decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_9,decoder_decoded_andMatrixInput_10,
    decoder_decoded_andMatrixInput_11};
  wire [12:0] _decoder_decoded_T_4 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_lo_2};
  wire  _decoder_decoded_T_5 = &_decoder_decoded_T_4;
  wire  decoder_decoded_andMatrixInput_9_2 = decoder_decoded_invInputs[28];
  wire [5:0] decoder_decoded_lo_3 = {decoder_decoded_andMatrixInput_7,decoder_decoded_andMatrixInput_8,
    decoder_decoded_andMatrixInput_9_2,decoder_decoded_andMatrixInput_9,decoder_decoded_andMatrixInput_10,
    decoder_decoded_andMatrixInput_11};
  wire [12:0] _decoder_decoded_T_6 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_lo_3};
  wire  _decoder_decoded_T_7 = &_decoder_decoded_T_6;
  wire  decoder_decoded_andMatrixInput_2_4 = io_inst[2];
  wire  decoder_decoded_andMatrixInput_5_3 = decoder_decoded_invInputs[6];
  wire  decoder_decoded_andMatrixInput_6_3 = decoder_decoded_invInputs[12];
  wire  decoder_decoded_andMatrixInput_7_3 = io_inst[13];
  wire  decoder_decoded_andMatrixInput_8_3 = decoder_decoded_invInputs[14];
  wire [8:0] _decoder_decoded_T_8 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_4,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_2,
    decoder_decoded_andMatrixInput_5_3,decoder_decoded_andMatrixInput_6_3,decoder_decoded_andMatrixInput_7_3,
    decoder_decoded_andMatrixInput_8_3};
  wire  _decoder_decoded_T_9 = &_decoder_decoded_T_8;
  wire [9:0] _decoder_decoded_T_10 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_4,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_2,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_5_3,decoder_decoded_andMatrixInput_6_3,
    decoder_decoded_andMatrixInput_7_3,decoder_decoded_andMatrixInput_8_3};
  wire  _decoder_decoded_T_11 = &_decoder_decoded_T_10;
  wire  decoder_decoded_andMatrixInput_5_5 = io_inst[5];
  wire [9:0] _decoder_decoded_T_12 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_4,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_2,
    decoder_decoded_andMatrixInput_5_5,decoder_decoded_andMatrixInput_5_3,decoder_decoded_andMatrixInput_6_3,
    decoder_decoded_andMatrixInput_7_3,decoder_decoded_andMatrixInput_8_3};
  wire  _decoder_decoded_T_13 = &_decoder_decoded_T_12;
  wire  decoder_decoded_andMatrixInput_9_5 = io_inst[27];
  wire  decoder_decoded_andMatrixInput_10_3 = io_inst[28];
  wire [6:0] decoder_decoded_lo_7 = {decoder_decoded_andMatrixInput_7,decoder_decoded_andMatrixInput_8,
    decoder_decoded_andMatrixInput_9_5,decoder_decoded_andMatrixInput_10_3,decoder_decoded_andMatrixInput_9,
    decoder_decoded_andMatrixInput_10,decoder_decoded_andMatrixInput_11};
  wire [13:0] _decoder_decoded_T_14 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_lo_7};
  wire  _decoder_decoded_T_15 = &_decoder_decoded_T_14;
  wire  decoder_decoded_andMatrixInput_13_1 = io_inst[29];
  wire [6:0] decoder_decoded_lo_8 = {decoder_decoded_andMatrixInput_8_3,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_9_2,
    decoder_decoded_andMatrixInput_13_1,decoder_decoded_andMatrixInput_10};
  wire [14:0] _decoder_decoded_T_16 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_6_3,
    decoder_decoded_lo_8};
  wire  _decoder_decoded_T_17 = &_decoder_decoded_T_16;
  wire  decoder_decoded_andMatrixInput_7_8 = decoder_decoded_invInputs[13];
  wire [14:0] _decoder_decoded_T_18 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_7_8,
    decoder_decoded_lo_8};
  wire  _decoder_decoded_T_19 = &_decoder_decoded_T_18;
  wire [6:0] decoder_decoded_lo_10 = {decoder_decoded_andMatrixInput_8_3,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_2,decoder_decoded_andMatrixInput_13_1,
    decoder_decoded_andMatrixInput_10,decoder_decoded_andMatrixInput_11};
  wire [14:0] _decoder_decoded_T_20 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_7_8,
    decoder_decoded_lo_10};
  wire  _decoder_decoded_T_21 = &_decoder_decoded_T_20;
  wire [7:0] decoder_decoded_lo_11 = {decoder_decoded_andMatrixInput_8_3,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_9_2,
    decoder_decoded_andMatrixInput_13_1,decoder_decoded_andMatrixInput_10,decoder_decoded_andMatrixInput_11};
  wire [15:0] _decoder_decoded_T_22 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_6_3,
    decoder_decoded_lo_11};
  wire  _decoder_decoded_T_23 = &_decoder_decoded_T_22;
  wire [7:0] decoder_decoded_lo_12 = {decoder_decoded_andMatrixInput_8_3,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_5,decoder_decoded_andMatrixInput_9_2,
    decoder_decoded_andMatrixInput_13_1,decoder_decoded_andMatrixInput_10,decoder_decoded_andMatrixInput_11};
  wire [15:0] _decoder_decoded_T_24 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_7_8,
    decoder_decoded_lo_12};
  wire  _decoder_decoded_T_25 = &_decoder_decoded_T_24;
  wire  decoder_decoded_andMatrixInput_7_12 = decoder_decoded_invInputs[20];
  wire  decoder_decoded_andMatrixInput_8_12 = decoder_decoded_invInputs[21];
  wire  decoder_decoded_andMatrixInput_9_11 = decoder_decoded_invInputs[22];
  wire  decoder_decoded_andMatrixInput_10_9 = decoder_decoded_invInputs[23];
  wire  decoder_decoded_andMatrixInput_11_9 = decoder_decoded_invInputs[24];
  wire  decoder_decoded_andMatrixInput_17 = io_inst[30];
  wire [9:0] decoder_decoded_hi_13 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_7_12,
    decoder_decoded_andMatrixInput_8_12,decoder_decoded_andMatrixInput_9_11};
  wire [18:0] _decoder_decoded_T_26 = {decoder_decoded_hi_13,decoder_decoded_andMatrixInput_10_9,
    decoder_decoded_andMatrixInput_11_9,decoder_decoded_andMatrixInput_7,decoder_decoded_andMatrixInput_8,
    decoder_decoded_andMatrixInput_9_5,decoder_decoded_andMatrixInput_10_3,decoder_decoded_andMatrixInput_9,
    decoder_decoded_andMatrixInput_17,decoder_decoded_andMatrixInput_11};
  wire  _decoder_decoded_T_27 = &_decoder_decoded_T_26;
  wire  decoder_decoded_andMatrixInput_15_3 = io_inst[31];
  wire [7:0] decoder_decoded_lo_14 = {decoder_decoded_andMatrixInput_8_3,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_9_2,
    decoder_decoded_andMatrixInput_13_1,decoder_decoded_andMatrixInput_10,decoder_decoded_andMatrixInput_15_3};
  wire [15:0] _decoder_decoded_T_28 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_6_3,
    decoder_decoded_lo_14};
  wire  _decoder_decoded_T_29 = &_decoder_decoded_T_28;
  wire [15:0] _decoder_decoded_T_30 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_7_8,
    decoder_decoded_lo_14};
  wire  _decoder_decoded_T_31 = &_decoder_decoded_T_30;
  wire [7:0] decoder_decoded_lo_16 = {decoder_decoded_andMatrixInput_10_9,decoder_decoded_andMatrixInput_11_9,
    decoder_decoded_andMatrixInput_7,decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_1,
    decoder_decoded_andMatrixInput_9,decoder_decoded_andMatrixInput_17,decoder_decoded_andMatrixInput_15_3};
  wire [15:0] _decoder_decoded_T_32 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_9_11,
    decoder_decoded_lo_16};
  wire  _decoder_decoded_T_33 = &_decoder_decoded_T_32;
  wire [7:0] decoder_decoded_lo_17 = {decoder_decoded_andMatrixInput_11_9,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_9_2,
    decoder_decoded_andMatrixInput_9,decoder_decoded_andMatrixInput_17,decoder_decoded_andMatrixInput_15_3};
  wire [16:0] _decoder_decoded_T_34 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_9_11,
    decoder_decoded_andMatrixInput_10_9,decoder_decoded_lo_17};
  wire  _decoder_decoded_T_35 = &_decoder_decoded_T_34;
  wire [7:0] decoder_decoded_lo_18 = {decoder_decoded_andMatrixInput_11_9,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_10_3,
    decoder_decoded_andMatrixInput_9,decoder_decoded_andMatrixInput_17,decoder_decoded_andMatrixInput_15_3};
  wire [16:0] _decoder_decoded_T_36 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_9_11,
    decoder_decoded_andMatrixInput_10_9,decoder_decoded_lo_18};
  wire  _decoder_decoded_T_37 = &_decoder_decoded_T_36;
  wire [9:0] decoder_decoded_lo_19 = {decoder_decoded_andMatrixInput_9_11,decoder_decoded_andMatrixInput_10_9,
    decoder_decoded_andMatrixInput_11_9,decoder_decoded_andMatrixInput_7,decoder_decoded_andMatrixInput_8,
    decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_9_2,decoder_decoded_andMatrixInput_13_1,
    decoder_decoded_andMatrixInput_17,decoder_decoded_andMatrixInput_15_3};
  wire [4:0] decoder_decoded_hi_lo_18 = {decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_7_8,
    decoder_decoded_andMatrixInput_8_3,decoder_decoded_andMatrixInput_7_12,decoder_decoded_andMatrixInput_8_12};
  wire [20:0] _decoder_decoded_T_38 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_hi_lo_18,decoder_decoded_lo_19};
  wire  _decoder_decoded_T_39 = &_decoder_decoded_T_38;
  wire [4:0] decoder_decoded_lo_lo_19 = {decoder_decoded_andMatrixInput_9_1,decoder_decoded_andMatrixInput_10_3,
    decoder_decoded_andMatrixInput_13_1,decoder_decoded_andMatrixInput_17,decoder_decoded_andMatrixInput_15_3};
  wire [10:0] decoder_decoded_lo_20 = {decoder_decoded_andMatrixInput_8_12,decoder_decoded_andMatrixInput_9_11,
    decoder_decoded_andMatrixInput_10_9,decoder_decoded_andMatrixInput_11_9,decoder_decoded_andMatrixInput_7,
    decoder_decoded_andMatrixInput_8,decoder_decoded_lo_lo_19};
  wire [4:0] decoder_decoded_hi_lo_19 = {decoder_decoded_andMatrixInput_4,decoder_decoded_andMatrixInput_6_3,
    decoder_decoded_andMatrixInput_7_8,decoder_decoded_andMatrixInput_8_3,decoder_decoded_andMatrixInput_7_12};
  wire [21:0] _decoder_decoded_T_40 = {decoder_decoded_andMatrixInput_0,decoder_decoded_andMatrixInput_1,
    decoder_decoded_andMatrixInput_2_1,decoder_decoded_andMatrixInput_3_1,decoder_decoded_andMatrixInput_4_1,
    decoder_decoded_andMatrixInput_3,decoder_decoded_hi_lo_19,decoder_decoded_lo_20};
  wire  _decoder_decoded_T_41 = &_decoder_decoded_T_40;
  wire [6:0] _decoder_decoded_orMatrixOutputs_T = {_decoder_decoded_T_1,_decoder_decoded_T_3,_decoder_decoded_T_25,
    _decoder_decoded_T_27,_decoder_decoded_T_29,_decoder_decoded_T_31,_decoder_decoded_T_33};
  wire  _decoder_decoded_orMatrixOutputs_T_1 = |_decoder_decoded_orMatrixOutputs_T;
  wire  _decoder_decoded_orMatrixOutputs_T_2 = |_decoder_decoded_T_27;
  wire  _decoder_decoded_orMatrixOutputs_T_3 = |_decoder_decoded_T_15;
  wire [2:0] _decoder_decoded_orMatrixOutputs_T_4 = {_decoder_decoded_T_1,_decoder_decoded_T_5,_decoder_decoded_T_7};
  wire  _decoder_decoded_orMatrixOutputs_T_5 = |_decoder_decoded_orMatrixOutputs_T_4;
  wire [1:0] _decoder_decoded_orMatrixOutputs_T_6 = {_decoder_decoded_T_21,_decoder_decoded_T_23};
  wire  _decoder_decoded_orMatrixOutputs_T_7 = |_decoder_decoded_orMatrixOutputs_T_6;
  wire [4:0] _decoder_decoded_orMatrixOutputs_T_8 = {_decoder_decoded_T_13,_decoder_decoded_T_29,_decoder_decoded_T_31,
    _decoder_decoded_T_35,_decoder_decoded_T_39};
  wire  _decoder_decoded_orMatrixOutputs_T_9 = |_decoder_decoded_orMatrixOutputs_T_8;
  wire [1:0] _decoder_decoded_orMatrixOutputs_T_10 = {_decoder_decoded_T_37,_decoder_decoded_T_41};
  wire  _decoder_decoded_orMatrixOutputs_T_11 = |_decoder_decoded_orMatrixOutputs_T_10;
  wire  _decoder_decoded_orMatrixOutputs_T_12 = |_decoder_decoded_T_7;
  wire  _decoder_decoded_orMatrixOutputs_T_13 = |_decoder_decoded_T_13;
  wire  _decoder_decoded_orMatrixOutputs_T_14 = |_decoder_decoded_T_1;
  wire [5:0] _decoder_decoded_orMatrixOutputs_T_15 = {_decoder_decoded_T_1,_decoder_decoded_T_3,_decoder_decoded_T_13,
    _decoder_decoded_T_17,_decoder_decoded_T_19,_decoder_decoded_T_21};
  wire  _decoder_decoded_orMatrixOutputs_T_16 = |_decoder_decoded_orMatrixOutputs_T_15;
  wire [7:0] _decoder_decoded_orMatrixOutputs_T_17 = {_decoder_decoded_T_1,_decoder_decoded_T_3,_decoder_decoded_T_17,
    _decoder_decoded_T_19,_decoder_decoded_T_21,_decoder_decoded_T_27,_decoder_decoded_T_35,_decoder_decoded_T_39};
  wire  _decoder_decoded_orMatrixOutputs_T_18 = |_decoder_decoded_orMatrixOutputs_T_17;
  wire [7:0] _decoder_decoded_orMatrixOutputs_T_19 = {_decoder_decoded_T_1,_decoder_decoded_T_3,_decoder_decoded_T_11,
    _decoder_decoded_T_21,_decoder_decoded_T_23,_decoder_decoded_T_27,_decoder_decoded_T_37,_decoder_decoded_T_41};
  wire  _decoder_decoded_orMatrixOutputs_T_20 = |_decoder_decoded_orMatrixOutputs_T_19;
  wire  _decoder_decoded_orMatrixOutputs_T_21 = |_decoder_decoded_T_9;
  wire [8:0] decoder_decoded_orMatrixOutputs_lo_5 = {2'h0,_decoder_decoded_orMatrixOutputs_T_11,
    _decoder_decoded_orMatrixOutputs_T_9,_decoder_decoded_orMatrixOutputs_T_7,_decoder_decoded_orMatrixOutputs_T_5,
    _decoder_decoded_orMatrixOutputs_T_3,_decoder_decoded_orMatrixOutputs_T_2,_decoder_decoded_orMatrixOutputs_T_1};
  wire [17:0] decoder_decoded_orMatrixOutputs = {_decoder_decoded_orMatrixOutputs_T_21,
    _decoder_decoded_orMatrixOutputs_T_20,_decoder_decoded_orMatrixOutputs_T_18,_decoder_decoded_orMatrixOutputs_T_16,
    _decoder_decoded_orMatrixOutputs_T_14,_decoder_decoded_orMatrixOutputs_T_13,_decoder_decoded_orMatrixOutputs_T_12,2'h0
    ,decoder_decoded_orMatrixOutputs_lo_5};
  wire [8:0] decoder_decoded_invMatrixOutputs_lo = {decoder_decoded_orMatrixOutputs[8],decoder_decoded_orMatrixOutputs[7
    ],decoder_decoded_orMatrixOutputs[6],decoder_decoded_orMatrixOutputs[5],decoder_decoded_orMatrixOutputs[4],
    decoder_decoded_orMatrixOutputs[3],decoder_decoded_orMatrixOutputs[2],decoder_decoded_orMatrixOutputs[1],
    decoder_decoded_orMatrixOutputs[0]};
  wire [17:0] decoder_decoded_invMatrixOutputs = {decoder_decoded_orMatrixOutputs[17],decoder_decoded_orMatrixOutputs[16
    ],decoder_decoded_orMatrixOutputs[15],decoder_decoded_orMatrixOutputs[14],decoder_decoded_orMatrixOutputs[13],
    decoder_decoded_orMatrixOutputs[12],decoder_decoded_orMatrixOutputs[11],decoder_decoded_orMatrixOutputs[10],
    decoder_decoded_orMatrixOutputs[9],decoder_decoded_invMatrixOutputs_lo};
  assign io_sigs_wen = decoder_decoded_invMatrixOutputs[16];
  assign io_sigs_ren1 = decoder_decoded_invMatrixOutputs[15];
  assign io_sigs_ren2 = decoder_decoded_invMatrixOutputs[14];
  assign io_sigs_ren3 = decoder_decoded_invMatrixOutputs[13];
  assign io_sigs_swap12 = decoder_decoded_invMatrixOutputs[12];
  assign io_sigs_swap23 = decoder_decoded_invMatrixOutputs[11];
  assign io_sigs_typeTagOut = decoder_decoded_invMatrixOutputs[8:7];
  assign io_sigs_fromint = decoder_decoded_invMatrixOutputs[6];
  assign io_sigs_toint = decoder_decoded_invMatrixOutputs[5];
  assign io_sigs_fastpipe = decoder_decoded_invMatrixOutputs[4];
  assign io_sigs_fma = decoder_decoded_invMatrixOutputs[3];
  assign io_sigs_div = decoder_decoded_invMatrixOutputs[2];
  assign io_sigs_sqrt = decoder_decoded_invMatrixOutputs[1];
  assign io_sigs_wflags = decoder_decoded_invMatrixOutputs[0];
endmodule