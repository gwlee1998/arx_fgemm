// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_393
`define RVX_GDEF_393

`define RVX_GDEF_422 6
`define RVX_GDEF_276 8
`define RVX_GDEF_411 3
`define RVX_GDEF_109 1

`define RVX_GDEF_302 (32'h 0)
`define RVX_GDEF_416 (32'h 8)
`define RVX_GDEF_271 (32'h 10)
`define RVX_GDEF_042 (32'h 18)
`define RVX_GDEF_237 (32'h 20)

`define RVX_GDEF_298 (`RVX_GDEF_302)
`define RVX_GDEF_198 (`RVX_GDEF_416)
`define RVX_GDEF_010 (`RVX_GDEF_271)
`define RVX_GDEF_097 (`RVX_GDEF_042)
`define RVX_GDEF_256 (`RVX_GDEF_237)

`define RVX_GDEF_334 5
`define RVX_GDEF_105 0
`define RVX_GDEF_342 9
`define RVX_GDEF_199 3
`define RVX_GDEF_139 7
`define RVX_GDEF_176 24

`define RVX_GDEF_136 32
`define RVX_GDEF_118 0

`define RVX_GDEF_106 32
`define RVX_GDEF_071 0

`define RVX_GDEF_243 32
`define RVX_GDEF_235 0

`define RVX_GDEF_048 32
`define RVX_GDEF_137 0

`endif