`ifndef __ERVP_CACHE_MEMORYMAP_OFFSET_H__
`define __ERVP_CACHE_MEMORYMAP_OFFSET_H__



// total
`define BW_MMAP_OFFSET_ERVP_CACHE 7
`define ERVP_CACHE_ADDR_INTERVAL 8
`define BW_UNUSED_ERVP_CACHE 3
`define NUM_ERVP_CACHE_SUBMODULE 1

// submodule cache
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START00 (32'h 0)
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START01 (32'h 8)
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START02 (32'h 10)
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START03 (32'h 18)
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST00 (32'h 20)
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST01 (32'h 28)
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST02 (32'h 30)
`define MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST03 (32'h 38)
`define MMAP_SUBOFFSET_CACHE_POLICY (32'h 40)
`define MMAP_SUBOFFSET_CACHE_BUSY (32'h 48)
`define MMAP_SUBOFFSET_CACHE_CONTROL_CMD (32'h 50)
`define MMAP_SUBOFFSET_CACHE_CONTROL_REGION_START (32'h 58)
`define MMAP_SUBOFFSET_CACHE_CONTROL_REGION_LAST (32'h 60)

`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_START00 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START00)
`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_START01 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START01)
`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_START02 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START02)
`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_START03 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_START03)
`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_LAST00 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST00)
`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_LAST01 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST01)
`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_LAST02 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST02)
`define MMAP_OFFSET_CACHE_CACHEABLE_REGION_LAST03 (`MMAP_SUBOFFSET_CACHE_CACHEABLE_REGION_LAST03)
`define MMAP_OFFSET_CACHE_POLICY (`MMAP_SUBOFFSET_CACHE_POLICY)
`define MMAP_OFFSET_CACHE_BUSY (`MMAP_SUBOFFSET_CACHE_BUSY)
`define MMAP_OFFSET_CACHE_CONTROL_CMD (`MMAP_SUBOFFSET_CACHE_CONTROL_CMD)
`define MMAP_OFFSET_CACHE_CONTROL_REGION_START (`MMAP_SUBOFFSET_CACHE_CONTROL_REGION_START)
`define MMAP_OFFSET_CACHE_CONTROL_REGION_LAST (`MMAP_SUBOFFSET_CACHE_CONTROL_REGION_LAST)

// reg cache.policy
`define BW_CACHE_POLICY 2
`define CACHE_POLICY_DEFAULT_VALUE 0
`define CACHE_POLICY_READ_ONLY 0
`define CACHE_POLICY_WRITE_THROUGH 1
`define CACHE_POLICY_WRITE_BACK 2
`define CACHE_POLICY_INDEX_WRITE_THROUGH 0
`define CACHE_POLICY_INDEX_WRITE_BACK 1

// reg cache.control_cmd
`define BW_CACHE_CONTROL_CMD 3
`define CACHE_CONTROL_CMD_DEFAULT_VALUE 0
`define CACHE_CONTROL_CMD_INITIALIZE 0
`define CACHE_CONTROL_CMD_INVALIDATE 1
`define CACHE_CONTROL_CMD_FLUSH 2
`define CACHE_CONTROL_CMD_CLEAN 3
`define CACHE_CONTROL_CMD_START 4
`define CACHE_CONTROL_CMD_STOP 5
`define CACHE_CONTROL_CMD_INDEX_INVALIDATE 0
`define CACHE_CONTROL_CMD_INDEX_FLUSH 1
`define CACHE_CONTROL_CMD_INDEX_START 2

// reg cache.cacheable_region_start
`define BW_CACHE_CACHEABLE_REGION_START 32
`define CACHE_CACHEABLE_REGION_START_DEFAULT_VALUE 0

// reg cache.cacheable_region_last
`define BW_CACHE_CACHEABLE_REGION_LAST 32
`define CACHE_CACHEABLE_REGION_LAST_DEFAULT_VALUE 0

// reg cache.busy
`define BW_CACHE_BUSY 1
`define CACHE_BUSY_DEFAULT_VALUE 0

// reg cache.control_region_start
`define BW_CACHE_CONTROL_REGION_START 32
`define CACHE_CONTROL_REGION_START_DEFAULT_VALUE 0

// reg cache.control_region_last
`define BW_CACHE_CONTROL_REGION_LAST 32
`define CACHE_CONTROL_REGION_LAST_DEFAULT_VALUE 0

`endif