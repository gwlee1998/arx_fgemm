`default_nettype wire
`include "timescale.vh"
module TLDebugModuleInner(
  input         clock,
  input         reset,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_opcode,
  input  [2:0]  auto_tl_in_a_bits_param,
  input  [1:0]  auto_tl_in_a_bits_size,
  input  [9:0]  auto_tl_in_a_bits_source,
  input  [11:0] auto_tl_in_a_bits_address,
  input  [3:0]  auto_tl_in_a_bits_mask,
  input  [31:0] auto_tl_in_a_bits_data,
  input         auto_tl_in_a_bits_corrupt,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_opcode,
  output [1:0]  auto_tl_in_d_bits_size,
  output [9:0]  auto_tl_in_d_bits_source,
  output [31:0] auto_tl_in_d_bits_data,
  output        auto_dmi_in_a_ready,
  input         auto_dmi_in_a_valid,
  input  [2:0]  auto_dmi_in_a_bits_opcode,
  input  [2:0]  auto_dmi_in_a_bits_param,
  input  [1:0]  auto_dmi_in_a_bits_size,
  input         auto_dmi_in_a_bits_source,
  input  [8:0]  auto_dmi_in_a_bits_address,
  input  [3:0]  auto_dmi_in_a_bits_mask,
  input  [31:0] auto_dmi_in_a_bits_data,
  input         auto_dmi_in_a_bits_corrupt,
  input         auto_dmi_in_d_ready,
  output        auto_dmi_in_d_valid,
  output [2:0]  auto_dmi_in_d_bits_opcode,
  output [1:0]  auto_dmi_in_d_bits_size,
  output        auto_dmi_in_d_bits_source,
  output [31:0] auto_dmi_in_d_bits_data,
  input         io_dmactive,
  output        io_innerCtrl_ready,
  input         io_innerCtrl_valid,
  input         io_innerCtrl_bits_resumereq,
  input  [9:0]  io_innerCtrl_bits_hartsel,
  input         io_innerCtrl_bits_ackhavereset,
  input         io_innerCtrl_bits_hrmask_0,
  output        io_hgDebugInt_0,
  input         io_hartIsInReset_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock;
  wire  monitor_reset;
  wire  monitor_io_in_a_ready;
  wire  monitor_io_in_a_valid;
  wire [2:0] monitor_io_in_a_bits_opcode;
  wire [2:0] monitor_io_in_a_bits_param;
  wire [1:0] monitor_io_in_a_bits_size;
  wire  monitor_io_in_a_bits_source;
  wire [8:0] monitor_io_in_a_bits_address;
  wire [3:0] monitor_io_in_a_bits_mask;
  wire  monitor_io_in_a_bits_corrupt;
  wire  monitor_io_in_d_ready;
  wire  monitor_io_in_d_valid;
  wire [2:0] monitor_io_in_d_bits_opcode;
  wire [1:0] monitor_io_in_d_bits_size;
  wire  monitor_io_in_d_bits_source;
  wire  monitor_1_clock;
  wire  monitor_1_reset;
  wire  monitor_1_io_in_a_ready;
  wire  monitor_1_io_in_a_valid;
  wire [2:0] monitor_1_io_in_a_bits_opcode;
  wire [2:0] monitor_1_io_in_a_bits_param;
  wire [1:0] monitor_1_io_in_a_bits_size;
  wire [9:0] monitor_1_io_in_a_bits_source;
  wire [11:0] monitor_1_io_in_a_bits_address;
  wire [3:0] monitor_1_io_in_a_bits_mask;
  wire  monitor_1_io_in_a_bits_corrupt;
  wire  monitor_1_io_in_d_ready;
  wire  monitor_1_io_in_d_valid;
  wire [2:0] monitor_1_io_in_d_bits_opcode;
  wire [1:0] monitor_1_io_in_d_bits_size;
  wire [9:0] monitor_1_io_in_d_bits_source;
  wire  hartIsInResetSync_0_debug_hartReset_0_clock;
  wire  hartIsInResetSync_0_debug_hartReset_0_reset;
  wire  hartIsInResetSync_0_debug_hartReset_0_io_d;
  wire  hartIsInResetSync_0_debug_hartReset_0_io_q;
  reg  haltedBitRegs;
  reg  resumeReqRegs;
  reg  haveResetBitRegs;
  wire  hamaskWrSel_0 = io_innerCtrl_bits_hartsel == 10'h0;
  reg  hrmaskReg_0;
  wire  _T_1 = ~io_dmactive;
  wire  _T_4 = io_innerCtrl_ready & io_innerCtrl_valid;
  reg  hrDebugIntReg_0;
  wire  _T_10 = ~haltedBitRegs;
  wire  _T_11 = hrDebugIntReg_0 & _T_10;
  wire  hartIsInResetSync_0 = hartIsInResetSync_0_debug_hartReset_0_io_q;
  wire  _T_12 = hartIsInResetSync_0 | _T_11;
  wire  _T_13 = hrmaskReg_0 & _T_12;
  wire  resumereq = _T_4 & io_innerCtrl_bits_resumereq;
  wire  _resumeAcks_T_1 = ~hamaskWrSel_0;
  wire  resumeAcks = resumereq ? ~resumeReqRegs & ~hamaskWrSel_0 : ~resumeReqRegs;
  wire [31:0] haltedStatus_0 = {{31'd0}, haltedBitRegs};
  wire  haltedSummary = |haltedStatus_0;
  wire [31:0] HALTSUM1RdData_haltsum1 = {{31'd0}, haltedSummary};
  reg [2:0] ABSTRACTCSReg_cmderr;
  wire  in_bits_read = auto_dmi_in_a_bits_opcode == 3'h4;
  wire [6:0] in_bits_index = auto_dmi_in_a_bits_address[8:2];
  wire [4:0] out_iindex = {in_bits_index[5],in_bits_index[3],in_bits_index[2],in_bits_index[1],in_bits_index[0]};
  wire [6:0] out_findex = in_bits_index & 7'h50;
  wire  _out_T_44 = out_findex == 7'h0;
  wire  _out_T_2 = out_findex == 7'h10;
  wire  _out_T_20 = out_findex == 7'h40;
  wire [31:0] _out_backSel_T = 32'h1 << out_iindex;
  wire  out_backSel_6 = _out_backSel_T[6];
  wire  out_woready__61 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_6 & out_findex == 7'h10
    ;
  wire [7:0] _out_backMask_T_11 = auto_dmi_in_a_bits_mask[3] ? 8'hff : 8'h0;
  wire [7:0] _out_backMask_T_9 = auto_dmi_in_a_bits_mask[2] ? 8'hff : 8'h0;
  wire [7:0] _out_backMask_T_7 = auto_dmi_in_a_bits_mask[1] ? 8'hff : 8'h0;
  wire [7:0] _out_backMask_T_5 = auto_dmi_in_a_bits_mask[0] ? 8'hff : 8'h0;
  wire [31:0] out_backMask = {_out_backMask_T_11,_out_backMask_T_9,_out_backMask_T_7,_out_backMask_T_5};
  wire  out_womask_61 = &out_backMask[10:8];
  wire  out_f_woready_61 = out_woready__61 & out_womask_61;
  reg [1:0] ctrlStateReg;
  wire  ABSTRACTCSWrEnLegal = ctrlStateReg == 2'h0;
  wire  ABSTRACTCSWrEn = out_f_woready_61 & ABSTRACTCSWrEnLegal;
  wire [2:0] ABSTRACTCSWrData_cmderr = auto_dmi_in_a_bits_data[10:8];
  wire [2:0] _ABSTRACTCSReg_cmderr_T = ~ABSTRACTCSWrData_cmderr;
  wire [2:0] _ABSTRACTCSReg_cmderr_T_1 = ABSTRACTCSReg_cmderr & _ABSTRACTCSReg_cmderr_T;
  wire [2:0] _GEN_37 = ABSTRACTCSWrEn ? _ABSTRACTCSReg_cmderr_T_1 : ABSTRACTCSReg_cmderr;
  wire  _T_1383 = ctrlStateReg == 2'h1;
  reg [7:0] COMMANDRdData_cmdtype;
  wire  commandRegIsAccessRegister = COMMANDRdData_cmdtype == 8'h0;
  reg [23:0] COMMANDRdData_control;
  wire [31:0] _accessRegisterCommandReg_T = {COMMANDRdData_cmdtype,COMMANDRdData_control};
  wire  accessRegisterCommandReg_transfer = _accessRegisterCommandReg_T[17];
  wire  accessRegisterCommandReg_write = _accessRegisterCommandReg_T[16];
  wire [15:0] accessRegisterCommandReg_regno = _accessRegisterCommandReg_T[15:0];
  wire [2:0] accessRegisterCommandReg_size = _accessRegisterCommandReg_T[22:20];
  wire  accessRegIsLegalSize = accessRegisterCommandReg_size == 3'h2 | accessRegisterCommandReg_size == 3'h3;
  wire  accessRegIsGPR = accessRegisterCommandReg_regno >= 16'h1000 & accessRegisterCommandReg_regno <= 16'h101f &
    accessRegIsLegalSize;
  wire  _GEN_3614 = ~accessRegisterCommandReg_transfer | accessRegIsGPR ? 1'h0 : 1'h1;
  wire  commandRegIsUnsupported = commandRegIsAccessRegister ? _GEN_3614 : 1'h1;
  wire  _GEN_3615 = (~accessRegisterCommandReg_transfer | accessRegIsGPR) & _T_10;
  wire  commandRegBadHaltResume = commandRegIsAccessRegister & _GEN_3615;
  wire  _GEN_3631 = commandRegIsUnsupported ? 1'h0 : commandRegBadHaltResume;
  wire  _GEN_3644 = ctrlStateReg == 2'h1 & _GEN_3631;
  wire  errorHaltResume = ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3644;
  wire [2:0] _GEN_38 = errorHaltResume ? 3'h4 : _GEN_37;
  wire  out_backSel_7 = _out_backSel_T[7];
  wire  out_woready__86 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_7 & out_findex == 7'h10
    ;
  wire  out_womask_86 = &out_backMask;
  wire  out_f_woready_86 = out_woready__86 & out_womask_86;
  wire  COMMANDWrEn = out_f_woready_86 & ABSTRACTCSWrEnLegal;
  wire [31:0] COMMANDWrDataVal = out_f_woready_86 ? auto_dmi_in_a_bits_data : 32'h0;
  wire [7:0] COMMANDWrData_cmdtype = COMMANDWrDataVal[31:24];
  wire  commandWrIsAccessRegister = COMMANDWrData_cmdtype == 8'h0;
  wire  _wrAccessRegisterCommand_T_1 = ABSTRACTCSReg_cmderr == 3'h0;
  wire  wrAccessRegisterCommand = COMMANDWrEn & commandWrIsAccessRegister & ABSTRACTCSReg_cmderr == 3'h0;
  wire  out_backSel_4 = _out_backSel_T[4];
  wire  out_woready__92 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_4 & out_findex == 7'h0
    ;
  wire  out_womask_92 = &out_backMask[7:0];
  wire  out_f_woready_92 = out_woready__92 & out_womask_92;
  wire  out_roready__92 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_4 & out_findex == 7'h0;
  wire  out_romask_92 = |out_backMask[7:0];
  wire  out_f_roready_92 = out_roready__92 & out_romask_92;
  wire  dmiAbstractDataAccessVec_0 = out_f_woready_92 | out_f_roready_92;
  reg [11:0] ABSTRACTAUTOReg_autoexecdata;
  wire  autoexecData_0 = dmiAbstractDataAccessVec_0 & ABSTRACTAUTOReg_autoexecdata[0];
  wire  out_backSel_16 = _out_backSel_T[16];
  wire  out_woready__27 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_16 & out_findex == 7'h0
    ;
  wire  out_f_woready_27 = out_woready__27 & out_womask_92;
  wire  out_roready__27 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_16 & out_findex == 7'h0
    ;
  wire  out_f_roready_27 = out_roready__27 & out_romask_92;
  wire  dmiProgramBufferAccessVec_0 = out_f_woready_27 | out_f_roready_27;
  reg [15:0] ABSTRACTAUTOReg_autoexecprogbuf;
  wire  autoexecProg_0 = dmiProgramBufferAccessVec_0 & ABSTRACTAUTOReg_autoexecprogbuf[0];
  wire  out_backSel_17 = _out_backSel_T[17];
  wire  out_woready__19 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_17 & out_findex == 7'h0
    ;
  wire  out_f_woready_19 = out_woready__19 & out_womask_92;
  wire  out_roready__19 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_17 & out_findex == 7'h0
    ;
  wire  out_f_roready_19 = out_roready__19 & out_romask_92;
  wire  dmiProgramBufferAccessVec_4 = out_f_woready_19 | out_f_roready_19;
  wire  autoexecProg_1 = dmiProgramBufferAccessVec_4 & ABSTRACTAUTOReg_autoexecprogbuf[1];
  wire  out_backSel_18 = _out_backSel_T[18];
  wire  out_woready__31 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_18 & out_findex == 7'h0
    ;
  wire  out_f_woready_31 = out_woready__31 & out_womask_92;
  wire  out_roready__31 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_18 & out_findex == 7'h0
    ;
  wire  out_f_roready_31 = out_roready__31 & out_romask_92;
  wire  dmiProgramBufferAccessVec_8 = out_f_woready_31 | out_f_roready_31;
  wire  autoexecProg_2 = dmiProgramBufferAccessVec_8 & ABSTRACTAUTOReg_autoexecprogbuf[2];
  wire  out_backSel_19 = _out_backSel_T[19];
  wire  out_woready__74 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_19 & out_findex == 7'h0
    ;
  wire  out_f_woready_74 = out_woready__74 & out_womask_92;
  wire  out_roready__74 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_19 & out_findex == 7'h0
    ;
  wire  out_f_roready_74 = out_roready__74 & out_romask_92;
  wire  dmiProgramBufferAccessVec_12 = out_f_woready_74 | out_f_roready_74;
  wire  autoexecProg_3 = dmiProgramBufferAccessVec_12 & ABSTRACTAUTOReg_autoexecprogbuf[3];
  wire  out_backSel_20 = _out_backSel_T[20];
  wire  out_woready__87 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_20 & out_findex == 7'h0
    ;
  wire  out_f_woready_87 = out_woready__87 & out_womask_92;
  wire  out_roready__87 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_20 & out_findex == 7'h0
    ;
  wire  out_f_roready_87 = out_roready__87 & out_romask_92;
  wire  dmiProgramBufferAccessVec_16 = out_f_woready_87 | out_f_roready_87;
  wire  autoexecProg_4 = dmiProgramBufferAccessVec_16 & ABSTRACTAUTOReg_autoexecprogbuf[4];
  wire  out_backSel_21 = _out_backSel_T[21];
  wire  out_woready__7 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_21 & out_findex == 7'h0
    ;
  wire  out_f_woready_7 = out_woready__7 & out_womask_92;
  wire  out_roready__7 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_21 & out_findex == 7'h0;
  wire  out_f_roready_7 = out_roready__7 & out_romask_92;
  wire  dmiProgramBufferAccessVec_20 = out_f_woready_7 | out_f_roready_7;
  wire  autoexecProg_5 = dmiProgramBufferAccessVec_20 & ABSTRACTAUTOReg_autoexecprogbuf[5];
  wire  out_backSel_22 = _out_backSel_T[22];
  wire  out_woready__15 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_22 & out_findex == 7'h0
    ;
  wire  out_f_woready_15 = out_woready__15 & out_womask_92;
  wire  out_roready__15 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_22 & out_findex == 7'h0
    ;
  wire  out_f_roready_15 = out_roready__15 & out_romask_92;
  wire  dmiProgramBufferAccessVec_24 = out_f_woready_15 | out_f_roready_15;
  wire  autoexecProg_6 = dmiProgramBufferAccessVec_24 & ABSTRACTAUTOReg_autoexecprogbuf[6];
  wire  out_backSel_23 = _out_backSel_T[23];
  wire  out_woready__70 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_23 & out_findex == 7'h0
    ;
  wire  out_f_woready_70 = out_woready__70 & out_womask_92;
  wire  out_roready__70 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_23 & out_findex == 7'h0
    ;
  wire  out_f_roready_70 = out_roready__70 & out_romask_92;
  wire  dmiProgramBufferAccessVec_28 = out_f_woready_70 | out_f_roready_70;
  wire  autoexecProg_7 = dmiProgramBufferAccessVec_28 & ABSTRACTAUTOReg_autoexecprogbuf[7];
  wire  out_backSel_24 = _out_backSel_T[24];
  wire  out_woready__82 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_24 & out_findex == 7'h0
    ;
  wire  out_f_woready_82 = out_woready__82 & out_womask_92;
  wire  out_roready__82 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_24 & out_findex == 7'h0
    ;
  wire  out_f_roready_82 = out_roready__82 & out_romask_92;
  wire  dmiProgramBufferAccessVec_32 = out_f_woready_82 | out_f_roready_82;
  wire  autoexecProg_8 = dmiProgramBufferAccessVec_32 & ABSTRACTAUTOReg_autoexecprogbuf[8];
  wire  out_backSel_25 = _out_backSel_T[25];
  wire  out_woready__23 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_25 & out_findex == 7'h0
    ;
  wire  out_f_woready_23 = out_woready__23 & out_womask_92;
  wire  out_roready__23 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_25 & out_findex == 7'h0
    ;
  wire  out_f_roready_23 = out_roready__23 & out_romask_92;
  wire  dmiProgramBufferAccessVec_36 = out_f_woready_23 | out_f_roready_23;
  wire  autoexecProg_9 = dmiProgramBufferAccessVec_36 & ABSTRACTAUTOReg_autoexecprogbuf[9];
  wire  out_backSel_26 = _out_backSel_T[26];
  wire  out_woready__0 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_26 & out_findex == 7'h0
    ;
  wire  out_f_woready = out_woready__0 & out_womask_92;
  wire  out_roready__0 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_26 & out_findex == 7'h0;
  wire  out_f_roready = out_roready__0 & out_romask_92;
  wire  dmiProgramBufferAccessVec_40 = out_f_woready | out_f_roready;
  wire  autoexecProg_10 = dmiProgramBufferAccessVec_40 & ABSTRACTAUTOReg_autoexecprogbuf[10];
  wire  out_backSel_27 = _out_backSel_T[27];
  wire  out_woready__78 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_27 & out_findex == 7'h0
    ;
  wire  out_f_woready_78 = out_woready__78 & out_womask_92;
  wire  out_roready__78 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_27 & out_findex == 7'h0
    ;
  wire  out_f_roready_78 = out_roready__78 & out_romask_92;
  wire  dmiProgramBufferAccessVec_44 = out_f_woready_78 | out_f_roready_78;
  wire  autoexecProg_11 = dmiProgramBufferAccessVec_44 & ABSTRACTAUTOReg_autoexecprogbuf[11];
  wire  out_backSel_28 = _out_backSel_T[28];
  wire  out_woready__66 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_28 & out_findex == 7'h0
    ;
  wire  out_f_woready_66 = out_woready__66 & out_womask_92;
  wire  out_roready__66 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_28 & out_findex == 7'h0
    ;
  wire  out_f_roready_66 = out_roready__66 & out_romask_92;
  wire  dmiProgramBufferAccessVec_48 = out_f_woready_66 | out_f_roready_66;
  wire  autoexecProg_12 = dmiProgramBufferAccessVec_48 & ABSTRACTAUTOReg_autoexecprogbuf[12];
  wire  out_backSel_29 = _out_backSel_T[29];
  wire  out_woready__35 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_29 & out_findex == 7'h0
    ;
  wire  out_f_woready_35 = out_woready__35 & out_womask_92;
  wire  out_roready__35 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_29 & out_findex == 7'h0
    ;
  wire  out_f_roready_35 = out_roready__35 & out_romask_92;
  wire  dmiProgramBufferAccessVec_52 = out_f_woready_35 | out_f_roready_35;
  wire  autoexecProg_13 = dmiProgramBufferAccessVec_52 & ABSTRACTAUTOReg_autoexecprogbuf[13];
  wire  out_backSel_30 = _out_backSel_T[30];
  wire  out_woready__11 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_30 & out_findex == 7'h0
    ;
  wire  out_f_woready_11 = out_woready__11 & out_womask_92;
  wire  out_roready__11 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_30 & out_findex == 7'h0
    ;
  wire  out_f_roready_11 = out_roready__11 & out_romask_92;
  wire  dmiProgramBufferAccessVec_56 = out_f_woready_11 | out_f_roready_11;
  wire  autoexecProg_14 = dmiProgramBufferAccessVec_56 & ABSTRACTAUTOReg_autoexecprogbuf[14];
  wire  out_backSel_31 = _out_backSel_T[31];
  wire  out_woready__96 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_31 & out_findex == 7'h0
    ;
  wire  out_f_woready_96 = out_woready__96 & out_womask_92;
  wire  out_roready__96 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & in_bits_read & out_backSel_31 & out_findex == 7'h0
    ;
  wire  out_f_roready_96 = out_roready__96 & out_romask_92;
  wire  dmiProgramBufferAccessVec_60 = out_f_woready_96 | out_f_roready_96;
  wire  autoexecProg_15 = dmiProgramBufferAccessVec_60 & ABSTRACTAUTOReg_autoexecprogbuf[15];
  wire  autoexec = autoexecData_0 | (autoexecProg_0 | autoexecProg_1 | autoexecProg_2 | autoexecProg_3 | autoexecProg_4
     | autoexecProg_5 | autoexecProg_6 | autoexecProg_7 | autoexecProg_8 | autoexecProg_9 | autoexecProg_10 |
    autoexecProg_11 | autoexecProg_12 | autoexecProg_13 | autoexecProg_14 | autoexecProg_15);
  wire  regAccessRegisterCommand = autoexec & commandRegIsAccessRegister & _wrAccessRegisterCommand_T_1;
  wire  commandWrIsUnsupported = COMMANDWrEn & ~commandWrIsAccessRegister;
  wire  _T_1382 = autoexec & commandRegIsUnsupported;
  wire  _GEN_3621 = commandWrIsUnsupported | _T_1382;
  wire  _GEN_3623 = wrAccessRegisterCommand | regAccessRegisterCommand ? 1'h0 : _GEN_3621;
  wire  _GEN_3642 = ctrlStateReg == 2'h1 & commandRegIsUnsupported;
  wire  errorUnsupported = ABSTRACTCSWrEnLegal ? _GEN_3623 : _GEN_3642;
  wire  _T_1384 = ctrlStateReg == 2'h2;
  wire  in_1_bits_read = auto_tl_in_a_bits_opcode == 3'h4;
  wire [9:0] in_1_bits_index = auto_tl_in_a_bits_address[11:2];
  wire [8:0] out_iindex_1 = {in_1_bits_index[8],in_1_bits_index[7],in_1_bits_index[6],in_1_bits_index[5],in_1_bits_index
    [4],in_1_bits_index[3],in_1_bits_index[2],in_1_bits_index[1],in_1_bits_index[0]};
  wire [9:0] out_findex_1 = in_1_bits_index & 10'h200;
  wire  _out_T_1122 = out_findex_1 == 10'h0;
  wire  _out_T_1642 = out_findex_1 == 10'h200;
  wire [511:0] _out_backSel_T_1 = 512'h1 << out_iindex_1;
  wire  out_backSel_67 = _out_backSel_T_1[67];
  wire  out_woready_1_841 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_backSel_67 & out_findex_1
     == 10'h0;
  wire [7:0] _out_backMask_T_23 = auto_tl_in_a_bits_mask[3] ? 8'hff : 8'h0;
  wire [7:0] _out_backMask_T_21 = auto_tl_in_a_bits_mask[2] ? 8'hff : 8'h0;
  wire [7:0] _out_backMask_T_19 = auto_tl_in_a_bits_mask[1] ? 8'hff : 8'h0;
  wire [7:0] _out_backMask_T_17 = auto_tl_in_a_bits_mask[0] ? 8'hff : 8'h0;
  wire [31:0] out_backMask_1 = {_out_backMask_T_23,_out_backMask_T_21,_out_backMask_T_19,_out_backMask_T_17};
  wire  out_womask_941 = &out_backMask_1[9:0];
  wire  out_f_woready_941 = out_woready_1_841 & out_womask_941;
  wire  _GEN_3640 = ctrlStateReg == 2'h2 & out_f_woready_941;
  wire  _GEN_3646 = ctrlStateReg == 2'h1 ? 1'h0 : _GEN_3640;
  wire  errorException = ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3646;
  wire  _errorBusy_T = ~ABSTRACTCSWrEnLegal;
  wire  out_backSel_8 = _out_backSel_T[8];
  wire  out_woready__4 = auto_dmi_in_a_valid & auto_dmi_in_d_ready & ~in_bits_read & out_backSel_8 & out_findex == 7'h10
    ;
  wire  out_womask_4 = &out_backMask[0];
  wire  out_f_woready_4 = out_woready__4 & out_womask_4;
  wire  _errorBusy_T_3 = out_f_woready_4 & _errorBusy_T;
  wire  _errorBusy_T_4 = out_f_woready_61 & ~ABSTRACTCSWrEnLegal | _errorBusy_T_3;
  wire  out_womask_6 = &out_backMask[31:16];
  wire  out_f_woready_6 = out_woready__4 & out_womask_6;
  wire  _errorBusy_T_6 = out_f_woready_6 & _errorBusy_T;
  wire  _errorBusy_T_7 = _errorBusy_T_4 | _errorBusy_T_6;
  wire  _errorBusy_T_9 = out_f_woready_86 & _errorBusy_T;
  wire  _errorBusy_T_10 = _errorBusy_T_7 | _errorBusy_T_9;
  wire  out_womask_93 = &out_backMask[15:8];
  wire  out_f_woready_93 = out_woready__92 & out_womask_93;
  wire  out_romask_93 = |out_backMask[15:8];
  wire  out_f_roready_93 = out_roready__92 & out_romask_93;
  wire  dmiAbstractDataAccessVec_1 = out_f_woready_93 | out_f_roready_93;
  wire  out_womask_94 = &out_backMask[23:16];
  wire  out_f_woready_94 = out_woready__92 & out_womask_94;
  wire  out_romask_94 = |out_backMask[23:16];
  wire  out_f_roready_94 = out_roready__92 & out_romask_94;
  wire  dmiAbstractDataAccessVec_2 = out_f_woready_94 | out_f_roready_94;
  wire  out_womask_95 = &out_backMask[31:24];
  wire  out_f_woready_95 = out_woready__92 & out_womask_95;
  wire  out_romask_95 = |out_backMask[31:24];
  wire  out_f_roready_95 = out_roready__92 & out_romask_95;
  wire  dmiAbstractDataAccessVec_3 = out_f_woready_95 | out_f_roready_95;
  wire  dmiAbstractDataAccess = dmiAbstractDataAccessVec_0 | dmiAbstractDataAccessVec_1 | dmiAbstractDataAccessVec_2 |
    dmiAbstractDataAccessVec_3;
  wire  _errorBusy_T_12 = dmiAbstractDataAccess & _errorBusy_T;
  wire  _errorBusy_T_13 = _errorBusy_T_10 | _errorBusy_T_12;
  wire  out_f_woready_28 = out_woready__27 & out_womask_93;
  wire  out_f_roready_28 = out_roready__27 & out_romask_93;
  wire  dmiProgramBufferAccessVec_1 = out_f_woready_28 | out_f_roready_28;
  wire  out_f_woready_29 = out_woready__27 & out_womask_94;
  wire  out_f_roready_29 = out_roready__27 & out_romask_94;
  wire  dmiProgramBufferAccessVec_2 = out_f_woready_29 | out_f_roready_29;
  wire  out_f_woready_30 = out_woready__27 & out_womask_95;
  wire  out_f_roready_30 = out_roready__27 & out_romask_95;
  wire  dmiProgramBufferAccessVec_3 = out_f_woready_30 | out_f_roready_30;
  wire  out_f_woready_20 = out_woready__19 & out_womask_93;
  wire  out_f_roready_20 = out_roready__19 & out_romask_93;
  wire  dmiProgramBufferAccessVec_5 = out_f_woready_20 | out_f_roready_20;
  wire  out_f_woready_21 = out_woready__19 & out_womask_94;
  wire  out_f_roready_21 = out_roready__19 & out_romask_94;
  wire  dmiProgramBufferAccessVec_6 = out_f_woready_21 | out_f_roready_21;
  wire  out_f_woready_22 = out_woready__19 & out_womask_95;
  wire  out_f_roready_22 = out_roready__19 & out_romask_95;
  wire  dmiProgramBufferAccessVec_7 = out_f_woready_22 | out_f_roready_22;
  wire  out_f_woready_32 = out_woready__31 & out_womask_93;
  wire  out_f_roready_32 = out_roready__31 & out_romask_93;
  wire  dmiProgramBufferAccessVec_9 = out_f_woready_32 | out_f_roready_32;
  wire  out_f_woready_33 = out_woready__31 & out_womask_94;
  wire  out_f_roready_33 = out_roready__31 & out_romask_94;
  wire  dmiProgramBufferAccessVec_10 = out_f_woready_33 | out_f_roready_33;
  wire  out_f_woready_34 = out_woready__31 & out_womask_95;
  wire  out_f_roready_34 = out_roready__31 & out_romask_95;
  wire  dmiProgramBufferAccessVec_11 = out_f_woready_34 | out_f_roready_34;
  wire  out_f_woready_75 = out_woready__74 & out_womask_93;
  wire  out_f_roready_75 = out_roready__74 & out_romask_93;
  wire  dmiProgramBufferAccessVec_13 = out_f_woready_75 | out_f_roready_75;
  wire  out_f_woready_76 = out_woready__74 & out_womask_94;
  wire  out_f_roready_76 = out_roready__74 & out_romask_94;
  wire  dmiProgramBufferAccessVec_14 = out_f_woready_76 | out_f_roready_76;
  wire  out_f_woready_77 = out_woready__74 & out_womask_95;
  wire  out_f_roready_77 = out_roready__74 & out_romask_95;
  wire  dmiProgramBufferAccessVec_15 = out_f_woready_77 | out_f_roready_77;
  wire  out_f_woready_88 = out_woready__87 & out_womask_93;
  wire  out_f_roready_88 = out_roready__87 & out_romask_93;
  wire  dmiProgramBufferAccessVec_17 = out_f_woready_88 | out_f_roready_88;
  wire  out_f_woready_89 = out_woready__87 & out_womask_94;
  wire  out_f_roready_89 = out_roready__87 & out_romask_94;
  wire  dmiProgramBufferAccessVec_18 = out_f_woready_89 | out_f_roready_89;
  wire  out_f_woready_90 = out_woready__87 & out_womask_95;
  wire  out_f_roready_90 = out_roready__87 & out_romask_95;
  wire  dmiProgramBufferAccessVec_19 = out_f_woready_90 | out_f_roready_90;
  wire  out_f_woready_8 = out_woready__7 & out_womask_93;
  wire  out_f_roready_8 = out_roready__7 & out_romask_93;
  wire  dmiProgramBufferAccessVec_21 = out_f_woready_8 | out_f_roready_8;
  wire  out_f_woready_9 = out_woready__7 & out_womask_94;
  wire  out_f_roready_9 = out_roready__7 & out_romask_94;
  wire  dmiProgramBufferAccessVec_22 = out_f_woready_9 | out_f_roready_9;
  wire  out_f_woready_10 = out_woready__7 & out_womask_95;
  wire  out_f_roready_10 = out_roready__7 & out_romask_95;
  wire  dmiProgramBufferAccessVec_23 = out_f_woready_10 | out_f_roready_10;
  wire  out_f_woready_16 = out_woready__15 & out_womask_93;
  wire  out_f_roready_16 = out_roready__15 & out_romask_93;
  wire  dmiProgramBufferAccessVec_25 = out_f_woready_16 | out_f_roready_16;
  wire  out_f_woready_17 = out_woready__15 & out_womask_94;
  wire  out_f_roready_17 = out_roready__15 & out_romask_94;
  wire  dmiProgramBufferAccessVec_26 = out_f_woready_17 | out_f_roready_17;
  wire  out_f_woready_18 = out_woready__15 & out_womask_95;
  wire  out_f_roready_18 = out_roready__15 & out_romask_95;
  wire  dmiProgramBufferAccessVec_27 = out_f_woready_18 | out_f_roready_18;
  wire  out_f_woready_71 = out_woready__70 & out_womask_93;
  wire  out_f_roready_71 = out_roready__70 & out_romask_93;
  wire  dmiProgramBufferAccessVec_29 = out_f_woready_71 | out_f_roready_71;
  wire  out_f_woready_72 = out_woready__70 & out_womask_94;
  wire  out_f_roready_72 = out_roready__70 & out_romask_94;
  wire  dmiProgramBufferAccessVec_30 = out_f_woready_72 | out_f_roready_72;
  wire  _dmiProgramBufferAccess_T_29 = dmiProgramBufferAccessVec_0 | dmiProgramBufferAccessVec_1 |
    dmiProgramBufferAccessVec_2 | dmiProgramBufferAccessVec_3 | dmiProgramBufferAccessVec_4 |
    dmiProgramBufferAccessVec_5 | dmiProgramBufferAccessVec_6 | dmiProgramBufferAccessVec_7 |
    dmiProgramBufferAccessVec_8 | dmiProgramBufferAccessVec_9 | dmiProgramBufferAccessVec_10 |
    dmiProgramBufferAccessVec_11 | dmiProgramBufferAccessVec_12 | dmiProgramBufferAccessVec_13 |
    dmiProgramBufferAccessVec_14 | dmiProgramBufferAccessVec_15 | dmiProgramBufferAccessVec_16 |
    dmiProgramBufferAccessVec_17 | dmiProgramBufferAccessVec_18 | dmiProgramBufferAccessVec_19 |
    dmiProgramBufferAccessVec_20 | dmiProgramBufferAccessVec_21 | dmiProgramBufferAccessVec_22 |
    dmiProgramBufferAccessVec_23 | dmiProgramBufferAccessVec_24 | dmiProgramBufferAccessVec_25 |
    dmiProgramBufferAccessVec_26 | dmiProgramBufferAccessVec_27 | dmiProgramBufferAccessVec_28 |
    dmiProgramBufferAccessVec_29 | dmiProgramBufferAccessVec_30;
  wire  out_f_woready_73 = out_woready__70 & out_womask_95;
  wire  out_f_roready_73 = out_roready__70 & out_romask_95;
  wire  dmiProgramBufferAccessVec_31 = out_f_woready_73 | out_f_roready_73;
  wire  out_f_woready_83 = out_woready__82 & out_womask_93;
  wire  out_f_roready_83 = out_roready__82 & out_romask_93;
  wire  dmiProgramBufferAccessVec_33 = out_f_woready_83 | out_f_roready_83;
  wire  out_f_woready_84 = out_woready__82 & out_womask_94;
  wire  out_f_roready_84 = out_roready__82 & out_romask_94;
  wire  dmiProgramBufferAccessVec_34 = out_f_woready_84 | out_f_roready_84;
  wire  out_f_woready_85 = out_woready__82 & out_womask_95;
  wire  out_f_roready_85 = out_roready__82 & out_romask_95;
  wire  dmiProgramBufferAccessVec_35 = out_f_woready_85 | out_f_roready_85;
  wire  out_f_woready_24 = out_woready__23 & out_womask_93;
  wire  out_f_roready_24 = out_roready__23 & out_romask_93;
  wire  dmiProgramBufferAccessVec_37 = out_f_woready_24 | out_f_roready_24;
  wire  out_f_woready_25 = out_woready__23 & out_womask_94;
  wire  out_f_roready_25 = out_roready__23 & out_romask_94;
  wire  dmiProgramBufferAccessVec_38 = out_f_woready_25 | out_f_roready_25;
  wire  out_f_woready_26 = out_woready__23 & out_womask_95;
  wire  out_f_roready_26 = out_roready__23 & out_romask_95;
  wire  dmiProgramBufferAccessVec_39 = out_f_woready_26 | out_f_roready_26;
  wire  out_f_woready_1 = out_woready__0 & out_womask_93;
  wire  out_f_roready_1 = out_roready__0 & out_romask_93;
  wire  dmiProgramBufferAccessVec_41 = out_f_woready_1 | out_f_roready_1;
  wire  out_f_woready_2 = out_woready__0 & out_womask_94;
  wire  out_f_roready_2 = out_roready__0 & out_romask_94;
  wire  dmiProgramBufferAccessVec_42 = out_f_woready_2 | out_f_roready_2;
  wire  out_f_woready_3 = out_woready__0 & out_womask_95;
  wire  out_f_roready_3 = out_roready__0 & out_romask_95;
  wire  dmiProgramBufferAccessVec_43 = out_f_woready_3 | out_f_roready_3;
  wire  out_f_woready_79 = out_woready__78 & out_womask_93;
  wire  out_f_roready_79 = out_roready__78 & out_romask_93;
  wire  dmiProgramBufferAccessVec_45 = out_f_woready_79 | out_f_roready_79;
  wire  out_f_woready_80 = out_woready__78 & out_womask_94;
  wire  out_f_roready_80 = out_roready__78 & out_romask_94;
  wire  dmiProgramBufferAccessVec_46 = out_f_woready_80 | out_f_roready_80;
  wire  out_f_woready_81 = out_woready__78 & out_womask_95;
  wire  out_f_roready_81 = out_roready__78 & out_romask_95;
  wire  dmiProgramBufferAccessVec_47 = out_f_woready_81 | out_f_roready_81;
  wire  out_f_woready_67 = out_woready__66 & out_womask_93;
  wire  out_f_roready_67 = out_roready__66 & out_romask_93;
  wire  dmiProgramBufferAccessVec_49 = out_f_woready_67 | out_f_roready_67;
  wire  out_f_woready_68 = out_woready__66 & out_womask_94;
  wire  out_f_roready_68 = out_roready__66 & out_romask_94;
  wire  dmiProgramBufferAccessVec_50 = out_f_woready_68 | out_f_roready_68;
  wire  out_f_woready_69 = out_woready__66 & out_womask_95;
  wire  out_f_roready_69 = out_roready__66 & out_romask_95;
  wire  dmiProgramBufferAccessVec_51 = out_f_woready_69 | out_f_roready_69;
  wire  out_f_woready_36 = out_woready__35 & out_womask_93;
  wire  out_f_roready_36 = out_roready__35 & out_romask_93;
  wire  dmiProgramBufferAccessVec_53 = out_f_woready_36 | out_f_roready_36;
  wire  out_f_woready_37 = out_woready__35 & out_womask_94;
  wire  out_f_roready_37 = out_roready__35 & out_romask_94;
  wire  dmiProgramBufferAccessVec_54 = out_f_woready_37 | out_f_roready_37;
  wire  out_f_woready_38 = out_woready__35 & out_womask_95;
  wire  out_f_roready_38 = out_roready__35 & out_romask_95;
  wire  dmiProgramBufferAccessVec_55 = out_f_woready_38 | out_f_roready_38;
  wire  out_f_woready_12 = out_woready__11 & out_womask_93;
  wire  out_f_roready_12 = out_roready__11 & out_romask_93;
  wire  dmiProgramBufferAccessVec_57 = out_f_woready_12 | out_f_roready_12;
  wire  out_f_woready_13 = out_woready__11 & out_womask_94;
  wire  out_f_roready_13 = out_roready__11 & out_romask_94;
  wire  dmiProgramBufferAccessVec_58 = out_f_woready_13 | out_f_roready_13;
  wire  out_f_woready_14 = out_woready__11 & out_womask_95;
  wire  out_f_roready_14 = out_roready__11 & out_romask_95;
  wire  dmiProgramBufferAccessVec_59 = out_f_woready_14 | out_f_roready_14;
  wire  _dmiProgramBufferAccess_T_59 = _dmiProgramBufferAccess_T_29 | dmiProgramBufferAccessVec_31 |
    dmiProgramBufferAccessVec_32 | dmiProgramBufferAccessVec_33 | dmiProgramBufferAccessVec_34 |
    dmiProgramBufferAccessVec_35 | dmiProgramBufferAccessVec_36 | dmiProgramBufferAccessVec_37 |
    dmiProgramBufferAccessVec_38 | dmiProgramBufferAccessVec_39 | dmiProgramBufferAccessVec_40 |
    dmiProgramBufferAccessVec_41 | dmiProgramBufferAccessVec_42 | dmiProgramBufferAccessVec_43 |
    dmiProgramBufferAccessVec_44 | dmiProgramBufferAccessVec_45 | dmiProgramBufferAccessVec_46 |
    dmiProgramBufferAccessVec_47 | dmiProgramBufferAccessVec_48 | dmiProgramBufferAccessVec_49 |
    dmiProgramBufferAccessVec_50 | dmiProgramBufferAccessVec_51 | dmiProgramBufferAccessVec_52 |
    dmiProgramBufferAccessVec_53 | dmiProgramBufferAccessVec_54 | dmiProgramBufferAccessVec_55 |
    dmiProgramBufferAccessVec_56 | dmiProgramBufferAccessVec_57 | dmiProgramBufferAccessVec_58 |
    dmiProgramBufferAccessVec_59 | dmiProgramBufferAccessVec_60;
  wire  out_f_woready_97 = out_woready__96 & out_womask_93;
  wire  out_f_roready_97 = out_roready__96 & out_romask_93;
  wire  dmiProgramBufferAccessVec_61 = out_f_woready_97 | out_f_roready_97;
  wire  out_f_woready_98 = out_woready__96 & out_womask_94;
  wire  out_f_roready_98 = out_roready__96 & out_romask_94;
  wire  dmiProgramBufferAccessVec_62 = out_f_woready_98 | out_f_roready_98;
  wire  out_f_woready_99 = out_woready__96 & out_womask_95;
  wire  out_f_roready_99 = out_roready__96 & out_romask_95;
  wire  dmiProgramBufferAccessVec_63 = out_f_woready_99 | out_f_roready_99;
  wire  dmiProgramBufferAccess = _dmiProgramBufferAccess_T_59 | dmiProgramBufferAccessVec_61 |
    dmiProgramBufferAccessVec_62 | dmiProgramBufferAccessVec_63;
  wire  _errorBusy_T_15 = dmiProgramBufferAccess & _errorBusy_T;
  wire  errorBusy = _errorBusy_T_13 | _errorBusy_T_15;
  wire [15:0] ABSTRACTAUTOWrData_autoexecprogbuf = auto_dmi_in_a_bits_data[31:16];
  wire [11:0] ABSTRACTAUTOWrData_autoexecdata = {{11'd0}, auto_dmi_in_a_bits_data[0]};
  wire [11:0] _ABSTRACTAUTOReg_autoexecdata_T = ABSTRACTAUTOWrData_autoexecdata & 12'h1;
  wire [23:0] COMMANDWrData_control = COMMANDWrDataVal[23:0];
  reg [7:0] abstractDataMem_0;
  reg [7:0] abstractDataMem_1;
  reg [7:0] abstractDataMem_2;
  reg [7:0] abstractDataMem_3;
  reg [7:0] programBufferMem_0;
  reg [7:0] programBufferMem_1;
  reg [7:0] programBufferMem_2;
  reg [7:0] programBufferMem_3;
  reg [7:0] programBufferMem_4;
  reg [7:0] programBufferMem_5;
  reg [7:0] programBufferMem_6;
  reg [7:0] programBufferMem_7;
  reg [7:0] programBufferMem_8;
  reg [7:0] programBufferMem_9;
  reg [7:0] programBufferMem_10;
  reg [7:0] programBufferMem_11;
  reg [7:0] programBufferMem_12;
  reg [7:0] programBufferMem_13;
  reg [7:0] programBufferMem_14;
  reg [7:0] programBufferMem_15;
  reg [7:0] programBufferMem_16;
  reg [7:0] programBufferMem_17;
  reg [7:0] programBufferMem_18;
  reg [7:0] programBufferMem_19;
  reg [7:0] programBufferMem_20;
  reg [7:0] programBufferMem_21;
  reg [7:0] programBufferMem_22;
  reg [7:0] programBufferMem_23;
  reg [7:0] programBufferMem_24;
  reg [7:0] programBufferMem_25;
  reg [7:0] programBufferMem_26;
  reg [7:0] programBufferMem_27;
  reg [7:0] programBufferMem_28;
  reg [7:0] programBufferMem_29;
  reg [7:0] programBufferMem_30;
  reg [7:0] programBufferMem_31;
  reg [7:0] programBufferMem_32;
  reg [7:0] programBufferMem_33;
  reg [7:0] programBufferMem_34;
  reg [7:0] programBufferMem_35;
  reg [7:0] programBufferMem_36;
  reg [7:0] programBufferMem_37;
  reg [7:0] programBufferMem_38;
  reg [7:0] programBufferMem_39;
  reg [7:0] programBufferMem_40;
  reg [7:0] programBufferMem_41;
  reg [7:0] programBufferMem_42;
  reg [7:0] programBufferMem_43;
  reg [7:0] programBufferMem_44;
  reg [7:0] programBufferMem_45;
  reg [7:0] programBufferMem_46;
  reg [7:0] programBufferMem_47;
  reg [7:0] programBufferMem_48;
  reg [7:0] programBufferMem_49;
  reg [7:0] programBufferMem_50;
  reg [7:0] programBufferMem_51;
  reg [7:0] programBufferMem_52;
  reg [7:0] programBufferMem_53;
  reg [7:0] programBufferMem_54;
  reg [7:0] programBufferMem_55;
  reg [7:0] programBufferMem_56;
  reg [7:0] programBufferMem_57;
  reg [7:0] programBufferMem_58;
  reg [7:0] programBufferMem_59;
  reg [7:0] programBufferMem_60;
  reg [7:0] programBufferMem_61;
  reg [7:0] programBufferMem_62;
  reg [7:0] programBufferMem_63;
  wire  _resumeReqRegs_T = ~hartIsInResetSync_0;
  wire  _resumeReqRegs_T_1 = resumeReqRegs & ~hartIsInResetSync_0;
  wire [1:0] _GEN_3655 = {{1'd0}, haltedBitRegs};
  wire [1:0] _haltedBitRegs_T = _GEN_3655 | 2'h1;
  wire [1:0] _GEN_3656 = {{1'd0}, _resumeReqRegs_T};
  wire [1:0] _haltedBitRegs_T_2 = _haltedBitRegs_T & _GEN_3656;
  wire [1:0] _haltedBitRegs_T_4 = _GEN_3655 & 2'h2;
  wire [1:0] _haltedBitRegs_T_6 = _haltedBitRegs_T_4 & _GEN_3656;
  wire  _haltedBitRegs_T_8 = haltedBitRegs & _resumeReqRegs_T;
  wire  out_backSel_66 = _out_backSel_T_1[66];
  wire  out_woready_1_708 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_backSel_66 & out_findex_1
     == 10'h0;
  wire  out_f_woready_808 = out_woready_1_708 & out_womask_941;
  wire [1:0] _GEN_61 = out_f_woready_808 ? _haltedBitRegs_T_6 : {{1'd0}, _haltedBitRegs_T_8};
  wire  out_backSel_64 = _out_backSel_T_1[64];
  wire  out_woready_1_547 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_backSel_64 & out_findex_1
     == 10'h0;
  wire  out_f_woready_647 = out_woready_1_547 & out_womask_941;
  wire [1:0] _GEN_62 = out_f_woready_647 ? _haltedBitRegs_T_2 : _GEN_61;
  wire [1:0] _GEN_3659 = {{1'd0}, resumeReqRegs};
  wire [1:0] _resumeReqRegs_T_3 = _GEN_3659 & 2'h2;
  wire [1:0] _resumeReqRegs_T_5 = _resumeReqRegs_T_3 & _GEN_3656;
  wire [1:0] _GEN_63 = out_f_woready_808 ? _resumeReqRegs_T_5 : {{1'd0}, _resumeReqRegs_T_1};
  wire  _resumeReqRegs_T_8 = (resumeReqRegs | hamaskWrSel_0) & _resumeReqRegs_T;
  wire [1:0] _GEN_64 = resumereq ? {{1'd0}, _resumeReqRegs_T_8} : _GEN_63;
  wire [1:0] _GEN_65 = _T_1 ? 2'h0 : _GEN_62;
  wire [1:0] _GEN_66 = _T_1 ? 2'h0 : _GEN_64;
  wire [31:0] out_prepend_2 = {programBufferMem_43,programBufferMem_42,programBufferMem_41,programBufferMem_40};
  wire [1:0] out_prepend_3 = {1'h0,ABSTRACTAUTOReg_autoexecdata[0]};
  wire [15:0] _out_T_108 = {{14'd0}, out_prepend_3};
  wire [31:0] out_prepend_4 = {ABSTRACTAUTOReg_autoexecprogbuf,_out_T_108};
  wire [31:0] out_prepend_7 = {programBufferMem_23,programBufferMem_22,programBufferMem_21,programBufferMem_20};
  wire [31:0] out_prepend_10 = {programBufferMem_59,programBufferMem_58,programBufferMem_57,programBufferMem_56};
  wire [31:0] out_prepend_13 = {programBufferMem_27,programBufferMem_26,programBufferMem_25,programBufferMem_24};
  wire [31:0] out_prepend_16 = {programBufferMem_7,programBufferMem_6,programBufferMem_5,programBufferMem_4};
  wire [31:0] out_prepend_19 = {programBufferMem_39,programBufferMem_38,programBufferMem_37,programBufferMem_36};
  wire [31:0] out_prepend_22 = {programBufferMem_3,programBufferMem_2,programBufferMem_1,programBufferMem_0};
  wire [31:0] out_prepend_25 = {programBufferMem_11,programBufferMem_10,programBufferMem_9,programBufferMem_8};
  wire [31:0] out_prepend_28 = {programBufferMem_55,programBufferMem_54,programBufferMem_53,programBufferMem_52};
  wire [16:0] out_prepend_41 = {resumeAcks,1'h0,1'h0,1'h0,1'h0,_T_10,_T_10,haltedBitRegs,haltedBitRegs,8'ha2};
  wire [20:0] out_prepend_45 = {1'h0,haveResetBitRegs,haveResetBitRegs,resumeAcks,out_prepend_41};
  wire [21:0] _out_T_642 = {{1'd0}, out_prepend_45};
  wire [22:0] out_prepend_46 = {1'h0,_out_T_642};
  wire  abstractCommandBusy = ctrlStateReg != 2'h0;
  wire [13:0] out_prepend_51 = {1'h0,abstractCommandBusy,1'h0,ABSTRACTCSReg_cmderr,8'h1};
  wire [23:0] _out_T_707 = {{10'd0}, out_prepend_51};
  wire [28:0] out_prepend_52 = {5'h10,_out_T_707};
  wire [31:0] out_prepend_55 = {programBufferMem_51,programBufferMem_50,programBufferMem_49,programBufferMem_48};
  wire [31:0] out_prepend_58 = {programBufferMem_31,programBufferMem_30,programBufferMem_29,programBufferMem_28};
  wire [31:0] out_prepend_61 = {programBufferMem_15,programBufferMem_14,programBufferMem_13,programBufferMem_12};
  wire [31:0] out_prepend_64 = {programBufferMem_47,programBufferMem_46,programBufferMem_45,programBufferMem_44};
  wire [31:0] out_prepend_67 = {programBufferMem_35,programBufferMem_34,programBufferMem_33,programBufferMem_32};
  wire [31:0] out_prepend_70 = {programBufferMem_19,programBufferMem_18,programBufferMem_17,programBufferMem_16};
  wire [31:0] out_prepend_73 = {abstractDataMem_3,abstractDataMem_2,abstractDataMem_1,abstractDataMem_0};
  wire [31:0] out_prepend_76 = {programBufferMem_63,programBufferMem_62,programBufferMem_61,programBufferMem_60};
  wire  _GEN_266 = 5'h1 == out_iindex ? _out_T_2 : _out_T_20;
  wire  _GEN_268 = 5'h3 == out_iindex ? _out_T_2 : 5'h2 == out_iindex | _GEN_266;
  wire  _GEN_269 = 5'h4 == out_iindex ? _out_T_44 : _GEN_268;
  wire  _GEN_271 = 5'h6 == out_iindex ? _out_T_2 : 5'h5 == out_iindex | _GEN_269;
  wire  _GEN_272 = 5'h7 == out_iindex ? _out_T_2 : _GEN_271;
  wire  _GEN_273 = 5'h8 == out_iindex ? _out_T_2 : _GEN_272;
  wire  _GEN_281 = 5'h10 == out_iindex ? _out_T_44 : 5'hf == out_iindex | (5'he == out_iindex | (5'hd == out_iindex | (5'hc
     == out_iindex | (5'hb == out_iindex | (5'ha == out_iindex | (5'h9 == out_iindex | _GEN_273))))));
  wire  _GEN_282 = 5'h11 == out_iindex ? _out_T_44 : _GEN_281;
  wire  _GEN_283 = 5'h12 == out_iindex ? _out_T_44 : _GEN_282;
  wire  _GEN_284 = 5'h13 == out_iindex ? _out_T_44 : _GEN_283;
  wire  _GEN_285 = 5'h14 == out_iindex ? _out_T_44 : _GEN_284;
  wire  _GEN_286 = 5'h15 == out_iindex ? _out_T_44 : _GEN_285;
  wire  _GEN_287 = 5'h16 == out_iindex ? _out_T_44 : _GEN_286;
  wire  _GEN_288 = 5'h17 == out_iindex ? _out_T_44 : _GEN_287;
  wire  _GEN_289 = 5'h18 == out_iindex ? _out_T_44 : _GEN_288;
  wire  _GEN_290 = 5'h19 == out_iindex ? _out_T_44 : _GEN_289;
  wire  _GEN_291 = 5'h1a == out_iindex ? _out_T_44 : _GEN_290;
  wire  _GEN_292 = 5'h1b == out_iindex ? _out_T_44 : _GEN_291;
  wire  _GEN_293 = 5'h1c == out_iindex ? _out_T_44 : _GEN_292;
  wire  _GEN_294 = 5'h1d == out_iindex ? _out_T_44 : _GEN_293;
  wire  _GEN_295 = 5'h1e == out_iindex ? _out_T_44 : _GEN_294;
  wire  _GEN_296 = 5'h1f == out_iindex ? _out_T_44 : _GEN_295;
  wire [31:0] _out_out_bits_data_WIRE_1_1 = {{9'd0}, out_prepend_46};
  wire [31:0] _GEN_298 = 5'h1 == out_iindex ? _out_out_bits_data_WIRE_1_1 : haltedStatus_0;
  wire [31:0] _GEN_299 = 5'h2 == out_iindex ? 32'h0 : _GEN_298;
  wire [31:0] _GEN_300 = 5'h3 == out_iindex ? HALTSUM1RdData_haltsum1 : _GEN_299;
  wire [31:0] _GEN_301 = 5'h4 == out_iindex ? out_prepend_73 : _GEN_300;
  wire [31:0] _GEN_302 = 5'h5 == out_iindex ? 32'h0 : _GEN_301;
  wire [31:0] _out_out_bits_data_WIRE_1_6 = {{3'd0}, out_prepend_52};
  wire [31:0] _GEN_303 = 5'h6 == out_iindex ? _out_out_bits_data_WIRE_1_6 : _GEN_302;
  wire [31:0] _GEN_304 = 5'h7 == out_iindex ? _accessRegisterCommandReg_T : _GEN_303;
  wire [31:0] _GEN_305 = 5'h8 == out_iindex ? out_prepend_4 : _GEN_304;
  wire [31:0] _GEN_306 = 5'h9 == out_iindex ? 32'h0 : _GEN_305;
  wire [31:0] _GEN_307 = 5'ha == out_iindex ? 32'h0 : _GEN_306;
  wire [31:0] _GEN_308 = 5'hb == out_iindex ? 32'h0 : _GEN_307;
  wire [31:0] _GEN_309 = 5'hc == out_iindex ? 32'h0 : _GEN_308;
  wire [31:0] _GEN_310 = 5'hd == out_iindex ? 32'h0 : _GEN_309;
  wire [31:0] _GEN_311 = 5'he == out_iindex ? 32'h0 : _GEN_310;
  wire [31:0] _GEN_312 = 5'hf == out_iindex ? 32'h0 : _GEN_311;
  wire [31:0] _GEN_313 = 5'h10 == out_iindex ? out_prepend_22 : _GEN_312;
  wire [31:0] _GEN_314 = 5'h11 == out_iindex ? out_prepend_16 : _GEN_313;
  wire [31:0] _GEN_315 = 5'h12 == out_iindex ? out_prepend_25 : _GEN_314;
  wire [31:0] _GEN_316 = 5'h13 == out_iindex ? out_prepend_61 : _GEN_315;
  wire [31:0] _GEN_317 = 5'h14 == out_iindex ? out_prepend_70 : _GEN_316;
  wire [31:0] _GEN_318 = 5'h15 == out_iindex ? out_prepend_7 : _GEN_317;
  wire [31:0] _GEN_319 = 5'h16 == out_iindex ? out_prepend_13 : _GEN_318;
  wire [31:0] _GEN_320 = 5'h17 == out_iindex ? out_prepend_58 : _GEN_319;
  wire [31:0] _GEN_321 = 5'h18 == out_iindex ? out_prepend_67 : _GEN_320;
  wire [31:0] _GEN_322 = 5'h19 == out_iindex ? out_prepend_19 : _GEN_321;
  wire [31:0] _GEN_323 = 5'h1a == out_iindex ? out_prepend_2 : _GEN_322;
  wire [31:0] _GEN_324 = 5'h1b == out_iindex ? out_prepend_64 : _GEN_323;
  wire [31:0] _GEN_325 = 5'h1c == out_iindex ? out_prepend_55 : _GEN_324;
  wire [31:0] _GEN_326 = 5'h1d == out_iindex ? out_prepend_28 : _GEN_325;
  wire [31:0] _GEN_327 = 5'h1e == out_iindex ? out_prepend_10 : _GEN_326;
  wire [31:0] _GEN_328 = 5'h1f == out_iindex ? out_prepend_76 : _GEN_327;
  reg  goReg;
  wire [9:0] hartGoingId = auto_tl_in_a_bits_data[9:0];
  wire  _T_341 = ~reset;
  wire  _T_342 = ~(hartGoingId == 10'h0);
  wire  out_backSel_65 = _out_backSel_T_1[65];
  wire  out_woready_1_370 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_backSel_65 & out_findex_1
     == 10'h0;
  wire  out_f_woready_470 = out_woready_1_370 & out_womask_941;
  wire  _GEN_397 = out_f_woready_470 ? 1'h0 : goReg;
  wire  _GEN_3628 = commandRegBadHaltResume ? 1'h0 : 1'h1;
  wire  _GEN_3632 = commandRegIsUnsupported ? 1'h0 : _GEN_3628;
  wire  _GEN_3645 = ctrlStateReg == 2'h1 & _GEN_3632;
  wire  goAbstract = ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3645;
  wire  _GEN_398 = goAbstract | _GEN_397;
  wire  accessRegisterCommandReg_postexec = _accessRegisterCommandReg_T[18];
  reg [31:0] abstractGeneratedMem_0;
  reg [31:0] abstractGeneratedMem_1;
  wire [15:0] _abstractGeneratedMem_0_inst_rd_T = accessRegisterCommandReg_regno & 16'h1f;
  wire [4:0] abstractGeneratedMem_0_inst_rd = _abstractGeneratedMem_0_inst_rd_T[4:0];
  wire [31:0] _abstractGeneratedMem_0_T = {17'h7000,accessRegisterCommandReg_size,abstractGeneratedMem_0_inst_rd,7'h3};
  wire [31:0] _abstractGeneratedMem_0_T_1 = {7'h1c,abstractGeneratedMem_0_inst_rd,5'h0,accessRegisterCommandReg_size,5'h0
    ,7'h23};
  wire  out_wimask_100 = &out_backMask_1[7:0];
  wire  out_wimask_101 = &out_backMask_1[15:8];
  wire  out_wimask_102 = &out_backMask_1[23:16];
  wire [23:0] out_prepend_78 = {6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
  wire  out_wimask_103 = &out_backMask_1[31:24];
  wire [31:0] out_prepend_79 = {6'h0,resumeReqRegs,goReg,out_prepend_78};
  wire  out_frontSel_217 = _out_backSel_T_1[217];
  wire  out_wivalid_1_40 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_217 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_140 = out_wivalid_1_40 & out_wimask_100;
  wire  out_f_wivalid_141 = out_wivalid_1_40 & out_wimask_101;
  wire  out_f_wivalid_142 = out_wivalid_1_40 & out_wimask_102;
  wire  out_f_wivalid_143 = out_wivalid_1_40 & out_wimask_103;
  wire  out_frontSel_216 = _out_backSel_T_1[216];
  wire  out_wivalid_1_176 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_216 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_276 = out_wivalid_1_176 & out_wimask_100;
  wire  out_f_wivalid_277 = out_wivalid_1_176 & out_wimask_101;
  wire  out_f_wivalid_278 = out_wivalid_1_176 & out_wimask_102;
  wire  out_f_wivalid_279 = out_wivalid_1_176 & out_wimask_103;
  wire  out_frontSel_211 = _out_backSel_T_1[211];
  wire  out_wivalid_1_200 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_211 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_300 = out_wivalid_1_200 & out_wimask_100;
  wire  out_f_wivalid_301 = out_wivalid_1_200 & out_wimask_101;
  wire  out_f_wivalid_302 = out_wivalid_1_200 & out_wimask_102;
  wire  out_f_wivalid_303 = out_wivalid_1_200 & out_wimask_103;
  wire  out_frontSel_221 = _out_backSel_T_1[221];
  wire  out_wivalid_1_232 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_221 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_332 = out_wivalid_1_232 & out_wimask_100;
  wire  out_f_wivalid_333 = out_wivalid_1_232 & out_wimask_101;
  wire  out_f_wivalid_334 = out_wivalid_1_232 & out_wimask_102;
  wire  out_f_wivalid_335 = out_wivalid_1_232 & out_wimask_103;
  wire  out_frontSel_220 = _out_backSel_T_1[220];
  wire  out_wivalid_1_309 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_220 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_409 = out_wivalid_1_309 & out_wimask_100;
  wire  out_f_wivalid_410 = out_wivalid_1_309 & out_wimask_101;
  wire  out_f_wivalid_411 = out_wivalid_1_309 & out_wimask_102;
  wire  out_f_wivalid_412 = out_wivalid_1_309 & out_wimask_103;
  wire  out_frontSel_224 = _out_backSel_T_1[224];
  wire  out_wivalid_1_403 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_224 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_503 = out_wivalid_1_403 & out_wimask_100;
  wire  out_f_wivalid_504 = out_wivalid_1_403 & out_wimask_101;
  wire  out_f_wivalid_505 = out_wivalid_1_403 & out_wimask_102;
  wire  out_f_wivalid_506 = out_wivalid_1_403 & out_wimask_103;
  wire  out_frontSel_212 = _out_backSel_T_1[212];
  wire  out_wivalid_1_467 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_212 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_567 = out_wivalid_1_467 & out_wimask_100;
  wire  out_f_wivalid_568 = out_wivalid_1_467 & out_wimask_101;
  wire  out_f_wivalid_569 = out_wivalid_1_467 & out_wimask_102;
  wire  out_f_wivalid_570 = out_wivalid_1_467 & out_wimask_103;
  wire  out_frontSel_219 = _out_backSel_T_1[219];
  wire  out_wivalid_1_624 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_219 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_724 = out_wivalid_1_624 & out_wimask_100;
  wire  out_f_wivalid_725 = out_wivalid_1_624 & out_wimask_101;
  wire  out_f_wivalid_726 = out_wivalid_1_624 & out_wimask_102;
  wire  out_f_wivalid_727 = out_wivalid_1_624 & out_wimask_103;
  wire  out_frontSel_208 = _out_backSel_T_1[208];
  wire  out_wivalid_1_668 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_208 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_768 = out_wivalid_1_668 & out_wimask_100;
  wire  out_f_wivalid_769 = out_wivalid_1_668 & out_wimask_101;
  wire  out_f_wivalid_770 = out_wivalid_1_668 & out_wimask_102;
  wire  out_f_wivalid_771 = out_wivalid_1_668 & out_wimask_103;
  wire  out_frontSel_213 = _out_backSel_T_1[213];
  wire  out_wivalid_1_696 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_213 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_796 = out_wivalid_1_696 & out_wimask_100;
  wire  out_f_wivalid_797 = out_wivalid_1_696 & out_wimask_101;
  wire  out_f_wivalid_798 = out_wivalid_1_696 & out_wimask_102;
  wire  out_f_wivalid_799 = out_wivalid_1_696 & out_wimask_103;
  wire  out_frontSel_223 = _out_backSel_T_1[223];
  wire  out_wivalid_1_733 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_223 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_833 = out_wivalid_1_733 & out_wimask_100;
  wire  out_f_wivalid_834 = out_wivalid_1_733 & out_wimask_101;
  wire  out_f_wivalid_835 = out_wivalid_1_733 & out_wimask_102;
  wire  out_f_wivalid_836 = out_wivalid_1_733 & out_wimask_103;
  wire  out_frontSel_209 = _out_backSel_T_1[209];
  wire  out_wivalid_1_785 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_209 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_885 = out_wivalid_1_785 & out_wimask_100;
  wire  out_f_wivalid_886 = out_wivalid_1_785 & out_wimask_101;
  wire  out_f_wivalid_887 = out_wivalid_1_785 & out_wimask_102;
  wire  out_f_wivalid_888 = out_wivalid_1_785 & out_wimask_103;
  wire  out_frontSel_218 = _out_backSel_T_1[218];
  wire  out_wivalid_1_918 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_218 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_1018 = out_wivalid_1_918 & out_wimask_100;
  wire  out_f_wivalid_1019 = out_wivalid_1_918 & out_wimask_101;
  wire  out_f_wivalid_1020 = out_wivalid_1_918 & out_wimask_102;
  wire  out_f_wivalid_1021 = out_wivalid_1_918 & out_wimask_103;
  wire  out_frontSel_214 = _out_backSel_T_1[214];
  wire  out_wivalid_1_991 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_214 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_1091 = out_wivalid_1_991 & out_wimask_100;
  wire  out_f_wivalid_1092 = out_wivalid_1_991 & out_wimask_101;
  wire  out_f_wivalid_1093 = out_wivalid_1_991 & out_wimask_102;
  wire  out_f_wivalid_1094 = out_wivalid_1_991 & out_wimask_103;
  wire  out_frontSel_210 = _out_backSel_T_1[210];
  wire  out_wivalid_1_1043 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_210 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_1143 = out_wivalid_1_1043 & out_wimask_100;
  wire  out_f_wivalid_1144 = out_wivalid_1_1043 & out_wimask_101;
  wire  out_f_wivalid_1145 = out_wivalid_1_1043 & out_wimask_102;
  wire  out_f_wivalid_1146 = out_wivalid_1_1043 & out_wimask_103;
  wire  out_frontSel_215 = _out_backSel_T_1[215];
  wire  out_wivalid_1_1159 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_215 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_1259 = out_wivalid_1_1159 & out_wimask_100;
  wire  out_f_wivalid_1260 = out_wivalid_1_1159 & out_wimask_101;
  wire  out_f_wivalid_1261 = out_wivalid_1_1159 & out_wimask_102;
  wire  out_f_wivalid_1262 = out_wivalid_1_1159 & out_wimask_103;
  wire  out_frontSel_222 = _out_backSel_T_1[222];
  wire  out_wivalid_1_1167 = auto_tl_in_a_valid & auto_tl_in_d_ready & ~in_1_bits_read & out_frontSel_222 & out_findex_1
     == 10'h0;
  wire  out_f_wivalid_1267 = out_wivalid_1_1167 & out_wimask_100;
  wire  out_f_wivalid_1268 = out_wivalid_1_1167 & out_wimask_101;
  wire  out_f_wivalid_1269 = out_wivalid_1_1167 & out_wimask_102;
  wire  out_f_wivalid_1270 = out_wivalid_1_1167 & out_wimask_103;
  wire  _GEN_2523 = 9'h1 == out_iindex_1 ? _out_T_1642 : _out_T_1642;
  wire  _GEN_2524 = 9'h2 == out_iindex_1 ? _out_T_1642 : _GEN_2523;
  wire  _GEN_2525 = 9'h3 == out_iindex_1 ? _out_T_1642 : _GEN_2524;
  wire  _GEN_2526 = 9'h4 == out_iindex_1 ? _out_T_1642 : _GEN_2525;
  wire  _GEN_2527 = 9'h5 == out_iindex_1 ? _out_T_1642 : _GEN_2526;
  wire  _GEN_2528 = 9'h6 == out_iindex_1 ? _out_T_1642 : _GEN_2527;
  wire  _GEN_2529 = 9'h7 == out_iindex_1 ? _out_T_1642 : _GEN_2528;
  wire  _GEN_2530 = 9'h8 == out_iindex_1 ? _out_T_1642 : _GEN_2529;
  wire  _GEN_2531 = 9'h9 == out_iindex_1 ? _out_T_1642 : _GEN_2530;
  wire  _GEN_2532 = 9'ha == out_iindex_1 ? _out_T_1642 : _GEN_2531;
  wire  _GEN_2533 = 9'hb == out_iindex_1 ? _out_T_1642 : _GEN_2532;
  wire  _GEN_2534 = 9'hc == out_iindex_1 ? _out_T_1642 : _GEN_2533;
  wire  _GEN_2535 = 9'hd == out_iindex_1 ? _out_T_1642 : _GEN_2534;
  wire  _GEN_2536 = 9'he == out_iindex_1 ? _out_T_1642 : _GEN_2535;
  wire  _GEN_2537 = 9'hf == out_iindex_1 ? _out_T_1642 : _GEN_2536;
  wire  _GEN_2538 = 9'h10 == out_iindex_1 ? _out_T_1642 : _GEN_2537;
  wire  _GEN_2539 = 9'h11 == out_iindex_1 ? _out_T_1642 : _GEN_2538;
  wire  _GEN_2540 = 9'h12 == out_iindex_1 ? _out_T_1642 : _GEN_2539;
  wire  _GEN_2541 = 9'h13 == out_iindex_1 ? _out_T_1642 : _GEN_2540;
  wire  _GEN_2542 = 9'h14 == out_iindex_1 ? _out_T_1642 : _GEN_2541;
  wire  _GEN_2557 = 9'h23 == out_iindex_1 | (9'h22 == out_iindex_1 | (9'h21 == out_iindex_1 | (9'h20 == out_iindex_1 | (9'h1f
     == out_iindex_1 | (9'h1e == out_iindex_1 | (9'h1d == out_iindex_1 | (9'h1c == out_iindex_1 | (9'h1b == out_iindex_1
     | (9'h1a == out_iindex_1 | (9'h19 == out_iindex_1 | (9'h18 == out_iindex_1 | (9'h17 == out_iindex_1 | (9'h16 ==
    out_iindex_1 | (9'h15 == out_iindex_1 | _GEN_2542))))))))))))));
  wire  _GEN_2572 = 9'h32 == out_iindex_1 | (9'h31 == out_iindex_1 | (9'h30 == out_iindex_1 | (9'h2f == out_iindex_1 | (9'h2e
     == out_iindex_1 | (9'h2d == out_iindex_1 | (9'h2c == out_iindex_1 | (9'h2b == out_iindex_1 | (9'h2a == out_iindex_1
     | (9'h29 == out_iindex_1 | (9'h28 == out_iindex_1 | (9'h27 == out_iindex_1 | (9'h26 == out_iindex_1 | (9'h25 ==
    out_iindex_1 | (9'h24 == out_iindex_1 | _GEN_2557))))))))))))));
  wire  _GEN_2586 = 9'h40 == out_iindex_1 ? _out_T_1122 : 9'h3f == out_iindex_1 | (9'h3e == out_iindex_1 | (9'h3d ==
    out_iindex_1 | (9'h3c == out_iindex_1 | (9'h3b == out_iindex_1 | (9'h3a == out_iindex_1 | (9'h39 == out_iindex_1 | (9'h38
     == out_iindex_1 | (9'h37 == out_iindex_1 | (9'h36 == out_iindex_1 | (9'h35 == out_iindex_1 | (9'h34 == out_iindex_1
     | (9'h33 == out_iindex_1 | _GEN_2572))))))))))));
  wire  _GEN_2587 = 9'h41 == out_iindex_1 ? _out_T_1122 : _GEN_2586;
  wire  _GEN_2588 = 9'h42 == out_iindex_1 ? _out_T_1122 : _GEN_2587;
  wire  _GEN_2589 = 9'h43 == out_iindex_1 ? _out_T_1122 : _GEN_2588;
  wire  _GEN_2604 = 9'h52 == out_iindex_1 | (9'h51 == out_iindex_1 | (9'h50 == out_iindex_1 | (9'h4f == out_iindex_1 | (9'h4e
     == out_iindex_1 | (9'h4d == out_iindex_1 | (9'h4c == out_iindex_1 | (9'h4b == out_iindex_1 | (9'h4a == out_iindex_1
     | (9'h49 == out_iindex_1 | (9'h48 == out_iindex_1 | (9'h47 == out_iindex_1 | (9'h46 == out_iindex_1 | (9'h45 ==
    out_iindex_1 | (9'h44 == out_iindex_1 | _GEN_2589))))))))))))));
  wire  _GEN_2619 = 9'h61 == out_iindex_1 | (9'h60 == out_iindex_1 | (9'h5f == out_iindex_1 | (9'h5e == out_iindex_1 | (9'h5d
     == out_iindex_1 | (9'h5c == out_iindex_1 | (9'h5b == out_iindex_1 | (9'h5a == out_iindex_1 | (9'h59 == out_iindex_1
     | (9'h58 == out_iindex_1 | (9'h57 == out_iindex_1 | (9'h56 == out_iindex_1 | (9'h55 == out_iindex_1 | (9'h54 ==
    out_iindex_1 | (9'h53 == out_iindex_1 | _GEN_2604))))))))))))));
  wire  _GEN_2634 = 9'h70 == out_iindex_1 | (9'h6f == out_iindex_1 | (9'h6e == out_iindex_1 | (9'h6d == out_iindex_1 | (9'h6c
     == out_iindex_1 | (9'h6b == out_iindex_1 | (9'h6a == out_iindex_1 | (9'h69 == out_iindex_1 | (9'h68 == out_iindex_1
     | (9'h67 == out_iindex_1 | (9'h66 == out_iindex_1 | (9'h65 == out_iindex_1 | (9'h64 == out_iindex_1 | (9'h63 ==
    out_iindex_1 | (9'h62 == out_iindex_1 | _GEN_2619))))))))))))));
  wire  _GEN_2649 = 9'h7f == out_iindex_1 | (9'h7e == out_iindex_1 | (9'h7d == out_iindex_1 | (9'h7c == out_iindex_1 | (9'h7b
     == out_iindex_1 | (9'h7a == out_iindex_1 | (9'h79 == out_iindex_1 | (9'h78 == out_iindex_1 | (9'h77 == out_iindex_1
     | (9'h76 == out_iindex_1 | (9'h75 == out_iindex_1 | (9'h74 == out_iindex_1 | (9'h73 == out_iindex_1 | (9'h72 ==
    out_iindex_1 | (9'h71 == out_iindex_1 | _GEN_2634))))))))))))));
  wire  _GEN_2664 = 9'h8e == out_iindex_1 | (9'h8d == out_iindex_1 | (9'h8c == out_iindex_1 | (9'h8b == out_iindex_1 | (9'h8a
     == out_iindex_1 | (9'h89 == out_iindex_1 | (9'h88 == out_iindex_1 | (9'h87 == out_iindex_1 | (9'h86 == out_iindex_1
     | (9'h85 == out_iindex_1 | (9'h84 == out_iindex_1 | (9'h83 == out_iindex_1 | (9'h82 == out_iindex_1 | (9'h81 ==
    out_iindex_1 | (9'h80 == out_iindex_1 | _GEN_2649))))))))))))));
  wire  _GEN_2679 = 9'h9d == out_iindex_1 | (9'h9c == out_iindex_1 | (9'h9b == out_iindex_1 | (9'h9a == out_iindex_1 | (9'h99
     == out_iindex_1 | (9'h98 == out_iindex_1 | (9'h97 == out_iindex_1 | (9'h96 == out_iindex_1 | (9'h95 == out_iindex_1
     | (9'h94 == out_iindex_1 | (9'h93 == out_iindex_1 | (9'h92 == out_iindex_1 | (9'h91 == out_iindex_1 | (9'h90 ==
    out_iindex_1 | (9'h8f == out_iindex_1 | _GEN_2664))))))))))))));
  wire  _GEN_2694 = 9'hac == out_iindex_1 | (9'hab == out_iindex_1 | (9'haa == out_iindex_1 | (9'ha9 == out_iindex_1 | (9'ha8
     == out_iindex_1 | (9'ha7 == out_iindex_1 | (9'ha6 == out_iindex_1 | (9'ha5 == out_iindex_1 | (9'ha4 == out_iindex_1
     | (9'ha3 == out_iindex_1 | (9'ha2 == out_iindex_1 | (9'ha1 == out_iindex_1 | (9'ha0 == out_iindex_1 | (9'h9f ==
    out_iindex_1 | (9'h9e == out_iindex_1 | _GEN_2679))))))))))))));
  wire  _GEN_2709 = 9'hbb == out_iindex_1 | (9'hba == out_iindex_1 | (9'hb9 == out_iindex_1 | (9'hb8 == out_iindex_1 | (9'hb7
     == out_iindex_1 | (9'hb6 == out_iindex_1 | (9'hb5 == out_iindex_1 | (9'hb4 == out_iindex_1 | (9'hb3 == out_iindex_1
     | (9'hb2 == out_iindex_1 | (9'hb1 == out_iindex_1 | (9'hb0 == out_iindex_1 | (9'haf == out_iindex_1 | (9'hae ==
    out_iindex_1 | (9'had == out_iindex_1 | _GEN_2694))))))))))))));
  wire  _GEN_2714 = 9'hc0 == out_iindex_1 ? _out_T_1122 : 9'hbf == out_iindex_1 | (9'hbe == out_iindex_1 | (9'hbd ==
    out_iindex_1 | (9'hbc == out_iindex_1 | _GEN_2709)));
  wire  _GEN_2728 = 9'hce == out_iindex_1 ? _out_T_1122 : 9'hcd == out_iindex_1 | (9'hcc == out_iindex_1 | (9'hcb ==
    out_iindex_1 | (9'hca == out_iindex_1 | (9'hc9 == out_iindex_1 | (9'hc8 == out_iindex_1 | (9'hc7 == out_iindex_1 | (9'hc6
     == out_iindex_1 | (9'hc5 == out_iindex_1 | (9'hc4 == out_iindex_1 | (9'hc3 == out_iindex_1 | (9'hc2 == out_iindex_1
     | (9'hc1 == out_iindex_1 | _GEN_2714))))))))))));
  wire  _GEN_2729 = 9'hcf == out_iindex_1 ? _out_T_1122 : _GEN_2728;
  wire  _GEN_2730 = 9'hd0 == out_iindex_1 ? _out_T_1122 : _GEN_2729;
  wire  _GEN_2731 = 9'hd1 == out_iindex_1 ? _out_T_1122 : _GEN_2730;
  wire  _GEN_2732 = 9'hd2 == out_iindex_1 ? _out_T_1122 : _GEN_2731;
  wire  _GEN_2733 = 9'hd3 == out_iindex_1 ? _out_T_1122 : _GEN_2732;
  wire  _GEN_2734 = 9'hd4 == out_iindex_1 ? _out_T_1122 : _GEN_2733;
  wire  _GEN_2735 = 9'hd5 == out_iindex_1 ? _out_T_1122 : _GEN_2734;
  wire  _GEN_2736 = 9'hd6 == out_iindex_1 ? _out_T_1122 : _GEN_2735;
  wire  _GEN_2737 = 9'hd7 == out_iindex_1 ? _out_T_1122 : _GEN_2736;
  wire  _GEN_2738 = 9'hd8 == out_iindex_1 ? _out_T_1122 : _GEN_2737;
  wire  _GEN_2739 = 9'hd9 == out_iindex_1 ? _out_T_1122 : _GEN_2738;
  wire  _GEN_2740 = 9'hda == out_iindex_1 ? _out_T_1122 : _GEN_2739;
  wire  _GEN_2741 = 9'hdb == out_iindex_1 ? _out_T_1122 : _GEN_2740;
  wire  _GEN_2742 = 9'hdc == out_iindex_1 ? _out_T_1122 : _GEN_2741;
  wire  _GEN_2743 = 9'hdd == out_iindex_1 ? _out_T_1122 : _GEN_2742;
  wire  _GEN_2744 = 9'hde == out_iindex_1 ? _out_T_1122 : _GEN_2743;
  wire  _GEN_2745 = 9'hdf == out_iindex_1 ? _out_T_1122 : _GEN_2744;
  wire  _GEN_2746 = 9'he0 == out_iindex_1 ? _out_T_1122 : _GEN_2745;
  wire  _GEN_2761 = 9'hef == out_iindex_1 | (9'hee == out_iindex_1 | (9'hed == out_iindex_1 | (9'hec == out_iindex_1 | (9'heb
     == out_iindex_1 | (9'hea == out_iindex_1 | (9'he9 == out_iindex_1 | (9'he8 == out_iindex_1 | (9'he7 == out_iindex_1
     | (9'he6 == out_iindex_1 | (9'he5 == out_iindex_1 | (9'he4 == out_iindex_1 | (9'he3 == out_iindex_1 | (9'he2 ==
    out_iindex_1 | (9'he1 == out_iindex_1 | _GEN_2746))))))))))))));
  wire  _GEN_2776 = 9'hfe == out_iindex_1 | (9'hfd == out_iindex_1 | (9'hfc == out_iindex_1 | (9'hfb == out_iindex_1 | (9'hfa
     == out_iindex_1 | (9'hf9 == out_iindex_1 | (9'hf8 == out_iindex_1 | (9'hf7 == out_iindex_1 | (9'hf6 == out_iindex_1
     | (9'hf5 == out_iindex_1 | (9'hf4 == out_iindex_1 | (9'hf3 == out_iindex_1 | (9'hf2 == out_iindex_1 | (9'hf1 ==
    out_iindex_1 | (9'hf0 == out_iindex_1 | _GEN_2761))))))))))))));
  wire  _GEN_2778 = 9'h100 == out_iindex_1 ? _out_T_1122 : 9'hff == out_iindex_1 | _GEN_2776;
  wire  _GEN_2779 = 9'h101 == out_iindex_1 ? _out_T_1122 : _GEN_2778;
  wire  _GEN_2780 = 9'h102 == out_iindex_1 ? _out_T_1122 : _GEN_2779;
  wire  _GEN_2781 = 9'h103 == out_iindex_1 ? _out_T_1122 : _GEN_2780;
  wire  _GEN_2782 = 9'h104 == out_iindex_1 ? _out_T_1122 : _GEN_2781;
  wire  _GEN_2783 = 9'h105 == out_iindex_1 ? _out_T_1122 : _GEN_2782;
  wire  _GEN_2784 = 9'h106 == out_iindex_1 ? _out_T_1122 : _GEN_2783;
  wire  _GEN_2785 = 9'h107 == out_iindex_1 ? _out_T_1122 : _GEN_2784;
  wire  _GEN_2786 = 9'h108 == out_iindex_1 ? _out_T_1122 : _GEN_2785;
  wire  _GEN_2787 = 9'h109 == out_iindex_1 ? _out_T_1122 : _GEN_2786;
  wire  _GEN_2788 = 9'h10a == out_iindex_1 ? _out_T_1122 : _GEN_2787;
  wire  _GEN_2789 = 9'h10b == out_iindex_1 ? _out_T_1122 : _GEN_2788;
  wire  _GEN_2790 = 9'h10c == out_iindex_1 ? _out_T_1122 : _GEN_2789;
  wire  _GEN_2791 = 9'h10d == out_iindex_1 ? _out_T_1122 : _GEN_2790;
  wire  _GEN_2792 = 9'h10e == out_iindex_1 ? _out_T_1122 : _GEN_2791;
  wire  _GEN_2793 = 9'h10f == out_iindex_1 ? _out_T_1122 : _GEN_2792;
  wire  _GEN_2794 = 9'h110 == out_iindex_1 ? _out_T_1122 : _GEN_2793;
  wire  _GEN_2795 = 9'h111 == out_iindex_1 ? _out_T_1122 : _GEN_2794;
  wire  _GEN_2796 = 9'h112 == out_iindex_1 ? _out_T_1122 : _GEN_2795;
  wire  _GEN_2797 = 9'h113 == out_iindex_1 ? _out_T_1122 : _GEN_2796;
  wire  _GEN_2798 = 9'h114 == out_iindex_1 ? _out_T_1122 : _GEN_2797;
  wire  _GEN_2799 = 9'h115 == out_iindex_1 ? _out_T_1122 : _GEN_2798;
  wire  _GEN_2800 = 9'h116 == out_iindex_1 ? _out_T_1122 : _GEN_2799;
  wire  _GEN_2801 = 9'h117 == out_iindex_1 ? _out_T_1122 : _GEN_2800;
  wire  _GEN_2802 = 9'h118 == out_iindex_1 ? _out_T_1122 : _GEN_2801;
  wire  _GEN_2803 = 9'h119 == out_iindex_1 ? _out_T_1122 : _GEN_2802;
  wire  _GEN_2804 = 9'h11a == out_iindex_1 ? _out_T_1122 : _GEN_2803;
  wire  _GEN_2805 = 9'h11b == out_iindex_1 ? _out_T_1122 : _GEN_2804;
  wire  _GEN_2806 = 9'h11c == out_iindex_1 ? _out_T_1122 : _GEN_2805;
  wire  _GEN_2807 = 9'h11d == out_iindex_1 ? _out_T_1122 : _GEN_2806;
  wire  _GEN_2808 = 9'h11e == out_iindex_1 ? _out_T_1122 : _GEN_2807;
  wire  _GEN_2809 = 9'h11f == out_iindex_1 ? _out_T_1122 : _GEN_2808;
  wire  _GEN_2810 = 9'h120 == out_iindex_1 ? _out_T_1122 : _GEN_2809;
  wire  _GEN_2811 = 9'h121 == out_iindex_1 ? _out_T_1122 : _GEN_2810;
  wire  _GEN_2812 = 9'h122 == out_iindex_1 ? _out_T_1122 : _GEN_2811;
  wire  _GEN_2813 = 9'h123 == out_iindex_1 ? _out_T_1122 : _GEN_2812;
  wire  _GEN_2814 = 9'h124 == out_iindex_1 ? _out_T_1122 : _GEN_2813;
  wire  _GEN_2815 = 9'h125 == out_iindex_1 ? _out_T_1122 : _GEN_2814;
  wire  _GEN_2816 = 9'h126 == out_iindex_1 ? _out_T_1122 : _GEN_2815;
  wire  _GEN_2817 = 9'h127 == out_iindex_1 ? _out_T_1122 : _GEN_2816;
  wire  _GEN_2818 = 9'h128 == out_iindex_1 ? _out_T_1122 : _GEN_2817;
  wire  _GEN_2819 = 9'h129 == out_iindex_1 ? _out_T_1122 : _GEN_2818;
  wire  _GEN_2820 = 9'h12a == out_iindex_1 ? _out_T_1122 : _GEN_2819;
  wire  _GEN_2821 = 9'h12b == out_iindex_1 ? _out_T_1122 : _GEN_2820;
  wire  _GEN_2822 = 9'h12c == out_iindex_1 ? _out_T_1122 : _GEN_2821;
  wire  _GEN_2823 = 9'h12d == out_iindex_1 ? _out_T_1122 : _GEN_2822;
  wire  _GEN_2824 = 9'h12e == out_iindex_1 ? _out_T_1122 : _GEN_2823;
  wire  _GEN_2825 = 9'h12f == out_iindex_1 ? _out_T_1122 : _GEN_2824;
  wire  _GEN_2826 = 9'h130 == out_iindex_1 ? _out_T_1122 : _GEN_2825;
  wire  _GEN_2827 = 9'h131 == out_iindex_1 ? _out_T_1122 : _GEN_2826;
  wire  _GEN_2828 = 9'h132 == out_iindex_1 ? _out_T_1122 : _GEN_2827;
  wire  _GEN_2829 = 9'h133 == out_iindex_1 ? _out_T_1122 : _GEN_2828;
  wire  _GEN_2830 = 9'h134 == out_iindex_1 ? _out_T_1122 : _GEN_2829;
  wire  _GEN_2831 = 9'h135 == out_iindex_1 ? _out_T_1122 : _GEN_2830;
  wire  _GEN_2832 = 9'h136 == out_iindex_1 ? _out_T_1122 : _GEN_2831;
  wire  _GEN_2833 = 9'h137 == out_iindex_1 ? _out_T_1122 : _GEN_2832;
  wire  _GEN_2834 = 9'h138 == out_iindex_1 ? _out_T_1122 : _GEN_2833;
  wire  _GEN_2835 = 9'h139 == out_iindex_1 ? _out_T_1122 : _GEN_2834;
  wire  _GEN_2836 = 9'h13a == out_iindex_1 ? _out_T_1122 : _GEN_2835;
  wire  _GEN_2837 = 9'h13b == out_iindex_1 ? _out_T_1122 : _GEN_2836;
  wire  _GEN_2838 = 9'h13c == out_iindex_1 ? _out_T_1122 : _GEN_2837;
  wire  _GEN_2839 = 9'h13d == out_iindex_1 ? _out_T_1122 : _GEN_2838;
  wire  _GEN_2840 = 9'h13e == out_iindex_1 ? _out_T_1122 : _GEN_2839;
  wire  _GEN_2841 = 9'h13f == out_iindex_1 ? _out_T_1122 : _GEN_2840;
  wire  _GEN_2842 = 9'h140 == out_iindex_1 ? _out_T_1122 : _GEN_2841;
  wire  _GEN_2843 = 9'h141 == out_iindex_1 ? _out_T_1122 : _GEN_2842;
  wire  _GEN_2844 = 9'h142 == out_iindex_1 ? _out_T_1122 : _GEN_2843;
  wire  _GEN_2845 = 9'h143 == out_iindex_1 ? _out_T_1122 : _GEN_2844;
  wire  _GEN_2846 = 9'h144 == out_iindex_1 ? _out_T_1122 : _GEN_2845;
  wire  _GEN_2847 = 9'h145 == out_iindex_1 ? _out_T_1122 : _GEN_2846;
  wire  _GEN_2848 = 9'h146 == out_iindex_1 ? _out_T_1122 : _GEN_2847;
  wire  _GEN_2849 = 9'h147 == out_iindex_1 ? _out_T_1122 : _GEN_2848;
  wire  _GEN_2850 = 9'h148 == out_iindex_1 ? _out_T_1122 : _GEN_2849;
  wire  _GEN_2851 = 9'h149 == out_iindex_1 ? _out_T_1122 : _GEN_2850;
  wire  _GEN_2852 = 9'h14a == out_iindex_1 ? _out_T_1122 : _GEN_2851;
  wire  _GEN_2853 = 9'h14b == out_iindex_1 ? _out_T_1122 : _GEN_2852;
  wire  _GEN_2854 = 9'h14c == out_iindex_1 ? _out_T_1122 : _GEN_2853;
  wire  _GEN_2855 = 9'h14d == out_iindex_1 ? _out_T_1122 : _GEN_2854;
  wire  _GEN_2856 = 9'h14e == out_iindex_1 ? _out_T_1122 : _GEN_2855;
  wire  _GEN_2857 = 9'h14f == out_iindex_1 ? _out_T_1122 : _GEN_2856;
  wire  _GEN_2858 = 9'h150 == out_iindex_1 ? _out_T_1122 : _GEN_2857;
  wire  _GEN_2859 = 9'h151 == out_iindex_1 ? _out_T_1122 : _GEN_2858;
  wire  _GEN_2860 = 9'h152 == out_iindex_1 ? _out_T_1122 : _GEN_2859;
  wire  _GEN_2861 = 9'h153 == out_iindex_1 ? _out_T_1122 : _GEN_2860;
  wire  _GEN_2862 = 9'h154 == out_iindex_1 ? _out_T_1122 : _GEN_2861;
  wire  _GEN_2863 = 9'h155 == out_iindex_1 ? _out_T_1122 : _GEN_2862;
  wire  _GEN_2864 = 9'h156 == out_iindex_1 ? _out_T_1122 : _GEN_2863;
  wire  _GEN_2865 = 9'h157 == out_iindex_1 ? _out_T_1122 : _GEN_2864;
  wire  _GEN_2866 = 9'h158 == out_iindex_1 ? _out_T_1122 : _GEN_2865;
  wire  _GEN_2867 = 9'h159 == out_iindex_1 ? _out_T_1122 : _GEN_2866;
  wire  _GEN_2868 = 9'h15a == out_iindex_1 ? _out_T_1122 : _GEN_2867;
  wire  _GEN_2869 = 9'h15b == out_iindex_1 ? _out_T_1122 : _GEN_2868;
  wire  _GEN_2870 = 9'h15c == out_iindex_1 ? _out_T_1122 : _GEN_2869;
  wire  _GEN_2871 = 9'h15d == out_iindex_1 ? _out_T_1122 : _GEN_2870;
  wire  _GEN_2872 = 9'h15e == out_iindex_1 ? _out_T_1122 : _GEN_2871;
  wire  _GEN_2873 = 9'h15f == out_iindex_1 ? _out_T_1122 : _GEN_2872;
  wire  _GEN_2874 = 9'h160 == out_iindex_1 ? _out_T_1122 : _GEN_2873;
  wire  _GEN_2875 = 9'h161 == out_iindex_1 ? _out_T_1122 : _GEN_2874;
  wire  _GEN_2876 = 9'h162 == out_iindex_1 ? _out_T_1122 : _GEN_2875;
  wire  _GEN_2877 = 9'h163 == out_iindex_1 ? _out_T_1122 : _GEN_2876;
  wire  _GEN_2878 = 9'h164 == out_iindex_1 ? _out_T_1122 : _GEN_2877;
  wire  _GEN_2879 = 9'h165 == out_iindex_1 ? _out_T_1122 : _GEN_2878;
  wire  _GEN_2880 = 9'h166 == out_iindex_1 ? _out_T_1122 : _GEN_2879;
  wire  _GEN_2881 = 9'h167 == out_iindex_1 ? _out_T_1122 : _GEN_2880;
  wire  _GEN_2882 = 9'h168 == out_iindex_1 ? _out_T_1122 : _GEN_2881;
  wire  _GEN_2883 = 9'h169 == out_iindex_1 ? _out_T_1122 : _GEN_2882;
  wire  _GEN_2884 = 9'h16a == out_iindex_1 ? _out_T_1122 : _GEN_2883;
  wire  _GEN_2885 = 9'h16b == out_iindex_1 ? _out_T_1122 : _GEN_2884;
  wire  _GEN_2886 = 9'h16c == out_iindex_1 ? _out_T_1122 : _GEN_2885;
  wire  _GEN_2887 = 9'h16d == out_iindex_1 ? _out_T_1122 : _GEN_2886;
  wire  _GEN_2888 = 9'h16e == out_iindex_1 ? _out_T_1122 : _GEN_2887;
  wire  _GEN_2889 = 9'h16f == out_iindex_1 ? _out_T_1122 : _GEN_2888;
  wire  _GEN_2890 = 9'h170 == out_iindex_1 ? _out_T_1122 : _GEN_2889;
  wire  _GEN_2891 = 9'h171 == out_iindex_1 ? _out_T_1122 : _GEN_2890;
  wire  _GEN_2892 = 9'h172 == out_iindex_1 ? _out_T_1122 : _GEN_2891;
  wire  _GEN_2893 = 9'h173 == out_iindex_1 ? _out_T_1122 : _GEN_2892;
  wire  _GEN_2894 = 9'h174 == out_iindex_1 ? _out_T_1122 : _GEN_2893;
  wire  _GEN_2895 = 9'h175 == out_iindex_1 ? _out_T_1122 : _GEN_2894;
  wire  _GEN_2896 = 9'h176 == out_iindex_1 ? _out_T_1122 : _GEN_2895;
  wire  _GEN_2897 = 9'h177 == out_iindex_1 ? _out_T_1122 : _GEN_2896;
  wire  _GEN_2898 = 9'h178 == out_iindex_1 ? _out_T_1122 : _GEN_2897;
  wire  _GEN_2899 = 9'h179 == out_iindex_1 ? _out_T_1122 : _GEN_2898;
  wire  _GEN_2900 = 9'h17a == out_iindex_1 ? _out_T_1122 : _GEN_2899;
  wire  _GEN_2901 = 9'h17b == out_iindex_1 ? _out_T_1122 : _GEN_2900;
  wire  _GEN_2902 = 9'h17c == out_iindex_1 ? _out_T_1122 : _GEN_2901;
  wire  _GEN_2903 = 9'h17d == out_iindex_1 ? _out_T_1122 : _GEN_2902;
  wire  _GEN_2904 = 9'h17e == out_iindex_1 ? _out_T_1122 : _GEN_2903;
  wire  _GEN_2905 = 9'h17f == out_iindex_1 ? _out_T_1122 : _GEN_2904;
  wire  _GEN_2906 = 9'h180 == out_iindex_1 ? _out_T_1122 : _GEN_2905;
  wire  _GEN_2907 = 9'h181 == out_iindex_1 ? _out_T_1122 : _GEN_2906;
  wire  _GEN_2908 = 9'h182 == out_iindex_1 ? _out_T_1122 : _GEN_2907;
  wire  _GEN_2909 = 9'h183 == out_iindex_1 ? _out_T_1122 : _GEN_2908;
  wire  _GEN_2910 = 9'h184 == out_iindex_1 ? _out_T_1122 : _GEN_2909;
  wire  _GEN_2911 = 9'h185 == out_iindex_1 ? _out_T_1122 : _GEN_2910;
  wire  _GEN_2912 = 9'h186 == out_iindex_1 ? _out_T_1122 : _GEN_2911;
  wire  _GEN_2913 = 9'h187 == out_iindex_1 ? _out_T_1122 : _GEN_2912;
  wire  _GEN_2914 = 9'h188 == out_iindex_1 ? _out_T_1122 : _GEN_2913;
  wire  _GEN_2915 = 9'h189 == out_iindex_1 ? _out_T_1122 : _GEN_2914;
  wire  _GEN_2916 = 9'h18a == out_iindex_1 ? _out_T_1122 : _GEN_2915;
  wire  _GEN_2917 = 9'h18b == out_iindex_1 ? _out_T_1122 : _GEN_2916;
  wire  _GEN_2918 = 9'h18c == out_iindex_1 ? _out_T_1122 : _GEN_2917;
  wire  _GEN_2919 = 9'h18d == out_iindex_1 ? _out_T_1122 : _GEN_2918;
  wire  _GEN_2920 = 9'h18e == out_iindex_1 ? _out_T_1122 : _GEN_2919;
  wire  _GEN_2921 = 9'h18f == out_iindex_1 ? _out_T_1122 : _GEN_2920;
  wire  _GEN_2922 = 9'h190 == out_iindex_1 ? _out_T_1122 : _GEN_2921;
  wire  _GEN_2923 = 9'h191 == out_iindex_1 ? _out_T_1122 : _GEN_2922;
  wire  _GEN_2924 = 9'h192 == out_iindex_1 ? _out_T_1122 : _GEN_2923;
  wire  _GEN_2925 = 9'h193 == out_iindex_1 ? _out_T_1122 : _GEN_2924;
  wire  _GEN_2926 = 9'h194 == out_iindex_1 ? _out_T_1122 : _GEN_2925;
  wire  _GEN_2927 = 9'h195 == out_iindex_1 ? _out_T_1122 : _GEN_2926;
  wire  _GEN_2928 = 9'h196 == out_iindex_1 ? _out_T_1122 : _GEN_2927;
  wire  _GEN_2929 = 9'h197 == out_iindex_1 ? _out_T_1122 : _GEN_2928;
  wire  _GEN_2930 = 9'h198 == out_iindex_1 ? _out_T_1122 : _GEN_2929;
  wire  _GEN_2931 = 9'h199 == out_iindex_1 ? _out_T_1122 : _GEN_2930;
  wire  _GEN_2932 = 9'h19a == out_iindex_1 ? _out_T_1122 : _GEN_2931;
  wire  _GEN_2933 = 9'h19b == out_iindex_1 ? _out_T_1122 : _GEN_2932;
  wire  _GEN_2934 = 9'h19c == out_iindex_1 ? _out_T_1122 : _GEN_2933;
  wire  _GEN_2935 = 9'h19d == out_iindex_1 ? _out_T_1122 : _GEN_2934;
  wire  _GEN_2936 = 9'h19e == out_iindex_1 ? _out_T_1122 : _GEN_2935;
  wire  _GEN_2937 = 9'h19f == out_iindex_1 ? _out_T_1122 : _GEN_2936;
  wire  _GEN_2938 = 9'h1a0 == out_iindex_1 ? _out_T_1122 : _GEN_2937;
  wire  _GEN_2939 = 9'h1a1 == out_iindex_1 ? _out_T_1122 : _GEN_2938;
  wire  _GEN_2940 = 9'h1a2 == out_iindex_1 ? _out_T_1122 : _GEN_2939;
  wire  _GEN_2941 = 9'h1a3 == out_iindex_1 ? _out_T_1122 : _GEN_2940;
  wire  _GEN_2942 = 9'h1a4 == out_iindex_1 ? _out_T_1122 : _GEN_2941;
  wire  _GEN_2943 = 9'h1a5 == out_iindex_1 ? _out_T_1122 : _GEN_2942;
  wire  _GEN_2944 = 9'h1a6 == out_iindex_1 ? _out_T_1122 : _GEN_2943;
  wire  _GEN_2945 = 9'h1a7 == out_iindex_1 ? _out_T_1122 : _GEN_2944;
  wire  _GEN_2946 = 9'h1a8 == out_iindex_1 ? _out_T_1122 : _GEN_2945;
  wire  _GEN_2947 = 9'h1a9 == out_iindex_1 ? _out_T_1122 : _GEN_2946;
  wire  _GEN_2948 = 9'h1aa == out_iindex_1 ? _out_T_1122 : _GEN_2947;
  wire  _GEN_2949 = 9'h1ab == out_iindex_1 ? _out_T_1122 : _GEN_2948;
  wire  _GEN_2950 = 9'h1ac == out_iindex_1 ? _out_T_1122 : _GEN_2949;
  wire  _GEN_2951 = 9'h1ad == out_iindex_1 ? _out_T_1122 : _GEN_2950;
  wire  _GEN_2952 = 9'h1ae == out_iindex_1 ? _out_T_1122 : _GEN_2951;
  wire  _GEN_2953 = 9'h1af == out_iindex_1 ? _out_T_1122 : _GEN_2952;
  wire  _GEN_2954 = 9'h1b0 == out_iindex_1 ? _out_T_1122 : _GEN_2953;
  wire  _GEN_2955 = 9'h1b1 == out_iindex_1 ? _out_T_1122 : _GEN_2954;
  wire  _GEN_2956 = 9'h1b2 == out_iindex_1 ? _out_T_1122 : _GEN_2955;
  wire  _GEN_2957 = 9'h1b3 == out_iindex_1 ? _out_T_1122 : _GEN_2956;
  wire  _GEN_2958 = 9'h1b4 == out_iindex_1 ? _out_T_1122 : _GEN_2957;
  wire  _GEN_2959 = 9'h1b5 == out_iindex_1 ? _out_T_1122 : _GEN_2958;
  wire  _GEN_2960 = 9'h1b6 == out_iindex_1 ? _out_T_1122 : _GEN_2959;
  wire  _GEN_2961 = 9'h1b7 == out_iindex_1 ? _out_T_1122 : _GEN_2960;
  wire  _GEN_2962 = 9'h1b8 == out_iindex_1 ? _out_T_1122 : _GEN_2961;
  wire  _GEN_2963 = 9'h1b9 == out_iindex_1 ? _out_T_1122 : _GEN_2962;
  wire  _GEN_2964 = 9'h1ba == out_iindex_1 ? _out_T_1122 : _GEN_2963;
  wire  _GEN_2965 = 9'h1bb == out_iindex_1 ? _out_T_1122 : _GEN_2964;
  wire  _GEN_2966 = 9'h1bc == out_iindex_1 ? _out_T_1122 : _GEN_2965;
  wire  _GEN_2967 = 9'h1bd == out_iindex_1 ? _out_T_1122 : _GEN_2966;
  wire  _GEN_2968 = 9'h1be == out_iindex_1 ? _out_T_1122 : _GEN_2967;
  wire  _GEN_2969 = 9'h1bf == out_iindex_1 ? _out_T_1122 : _GEN_2968;
  wire  _GEN_2970 = 9'h1c0 == out_iindex_1 ? _out_T_1122 : _GEN_2969;
  wire  _GEN_2971 = 9'h1c1 == out_iindex_1 ? _out_T_1122 : _GEN_2970;
  wire  _GEN_2972 = 9'h1c2 == out_iindex_1 ? _out_T_1122 : _GEN_2971;
  wire  _GEN_2973 = 9'h1c3 == out_iindex_1 ? _out_T_1122 : _GEN_2972;
  wire  _GEN_2974 = 9'h1c4 == out_iindex_1 ? _out_T_1122 : _GEN_2973;
  wire  _GEN_2975 = 9'h1c5 == out_iindex_1 ? _out_T_1122 : _GEN_2974;
  wire  _GEN_2976 = 9'h1c6 == out_iindex_1 ? _out_T_1122 : _GEN_2975;
  wire  _GEN_2977 = 9'h1c7 == out_iindex_1 ? _out_T_1122 : _GEN_2976;
  wire  _GEN_2978 = 9'h1c8 == out_iindex_1 ? _out_T_1122 : _GEN_2977;
  wire  _GEN_2979 = 9'h1c9 == out_iindex_1 ? _out_T_1122 : _GEN_2978;
  wire  _GEN_2980 = 9'h1ca == out_iindex_1 ? _out_T_1122 : _GEN_2979;
  wire  _GEN_2981 = 9'h1cb == out_iindex_1 ? _out_T_1122 : _GEN_2980;
  wire  _GEN_2982 = 9'h1cc == out_iindex_1 ? _out_T_1122 : _GEN_2981;
  wire  _GEN_2983 = 9'h1cd == out_iindex_1 ? _out_T_1122 : _GEN_2982;
  wire  _GEN_2984 = 9'h1ce == out_iindex_1 ? _out_T_1122 : _GEN_2983;
  wire  _GEN_2985 = 9'h1cf == out_iindex_1 ? _out_T_1122 : _GEN_2984;
  wire  _GEN_2986 = 9'h1d0 == out_iindex_1 ? _out_T_1122 : _GEN_2985;
  wire  _GEN_2987 = 9'h1d1 == out_iindex_1 ? _out_T_1122 : _GEN_2986;
  wire  _GEN_2988 = 9'h1d2 == out_iindex_1 ? _out_T_1122 : _GEN_2987;
  wire  _GEN_2989 = 9'h1d3 == out_iindex_1 ? _out_T_1122 : _GEN_2988;
  wire  _GEN_2990 = 9'h1d4 == out_iindex_1 ? _out_T_1122 : _GEN_2989;
  wire  _GEN_2991 = 9'h1d5 == out_iindex_1 ? _out_T_1122 : _GEN_2990;
  wire  _GEN_2992 = 9'h1d6 == out_iindex_1 ? _out_T_1122 : _GEN_2991;
  wire  _GEN_2993 = 9'h1d7 == out_iindex_1 ? _out_T_1122 : _GEN_2992;
  wire  _GEN_2994 = 9'h1d8 == out_iindex_1 ? _out_T_1122 : _GEN_2993;
  wire  _GEN_2995 = 9'h1d9 == out_iindex_1 ? _out_T_1122 : _GEN_2994;
  wire  _GEN_2996 = 9'h1da == out_iindex_1 ? _out_T_1122 : _GEN_2995;
  wire  _GEN_2997 = 9'h1db == out_iindex_1 ? _out_T_1122 : _GEN_2996;
  wire  _GEN_2998 = 9'h1dc == out_iindex_1 ? _out_T_1122 : _GEN_2997;
  wire  _GEN_2999 = 9'h1dd == out_iindex_1 ? _out_T_1122 : _GEN_2998;
  wire  _GEN_3000 = 9'h1de == out_iindex_1 ? _out_T_1122 : _GEN_2999;
  wire  _GEN_3001 = 9'h1df == out_iindex_1 ? _out_T_1122 : _GEN_3000;
  wire  _GEN_3002 = 9'h1e0 == out_iindex_1 ? _out_T_1122 : _GEN_3001;
  wire  _GEN_3003 = 9'h1e1 == out_iindex_1 ? _out_T_1122 : _GEN_3002;
  wire  _GEN_3004 = 9'h1e2 == out_iindex_1 ? _out_T_1122 : _GEN_3003;
  wire  _GEN_3005 = 9'h1e3 == out_iindex_1 ? _out_T_1122 : _GEN_3004;
  wire  _GEN_3006 = 9'h1e4 == out_iindex_1 ? _out_T_1122 : _GEN_3005;
  wire  _GEN_3007 = 9'h1e5 == out_iindex_1 ? _out_T_1122 : _GEN_3006;
  wire  _GEN_3008 = 9'h1e6 == out_iindex_1 ? _out_T_1122 : _GEN_3007;
  wire  _GEN_3009 = 9'h1e7 == out_iindex_1 ? _out_T_1122 : _GEN_3008;
  wire  _GEN_3010 = 9'h1e8 == out_iindex_1 ? _out_T_1122 : _GEN_3009;
  wire  _GEN_3011 = 9'h1e9 == out_iindex_1 ? _out_T_1122 : _GEN_3010;
  wire  _GEN_3012 = 9'h1ea == out_iindex_1 ? _out_T_1122 : _GEN_3011;
  wire  _GEN_3013 = 9'h1eb == out_iindex_1 ? _out_T_1122 : _GEN_3012;
  wire  _GEN_3014 = 9'h1ec == out_iindex_1 ? _out_T_1122 : _GEN_3013;
  wire  _GEN_3015 = 9'h1ed == out_iindex_1 ? _out_T_1122 : _GEN_3014;
  wire  _GEN_3016 = 9'h1ee == out_iindex_1 ? _out_T_1122 : _GEN_3015;
  wire  _GEN_3017 = 9'h1ef == out_iindex_1 ? _out_T_1122 : _GEN_3016;
  wire  _GEN_3018 = 9'h1f0 == out_iindex_1 ? _out_T_1122 : _GEN_3017;
  wire  _GEN_3019 = 9'h1f1 == out_iindex_1 ? _out_T_1122 : _GEN_3018;
  wire  _GEN_3020 = 9'h1f2 == out_iindex_1 ? _out_T_1122 : _GEN_3019;
  wire  _GEN_3021 = 9'h1f3 == out_iindex_1 ? _out_T_1122 : _GEN_3020;
  wire  _GEN_3022 = 9'h1f4 == out_iindex_1 ? _out_T_1122 : _GEN_3021;
  wire  _GEN_3023 = 9'h1f5 == out_iindex_1 ? _out_T_1122 : _GEN_3022;
  wire  _GEN_3024 = 9'h1f6 == out_iindex_1 ? _out_T_1122 : _GEN_3023;
  wire  _GEN_3025 = 9'h1f7 == out_iindex_1 ? _out_T_1122 : _GEN_3024;
  wire  _GEN_3026 = 9'h1f8 == out_iindex_1 ? _out_T_1122 : _GEN_3025;
  wire  _GEN_3027 = 9'h1f9 == out_iindex_1 ? _out_T_1122 : _GEN_3026;
  wire  _GEN_3028 = 9'h1fa == out_iindex_1 ? _out_T_1122 : _GEN_3027;
  wire  _GEN_3029 = 9'h1fb == out_iindex_1 ? _out_T_1122 : _GEN_3028;
  wire  _GEN_3030 = 9'h1fc == out_iindex_1 ? _out_T_1122 : _GEN_3029;
  wire  _GEN_3031 = 9'h1fd == out_iindex_1 ? _out_T_1122 : _GEN_3030;
  wire  _GEN_3032 = 9'h1fe == out_iindex_1 ? _out_T_1122 : _GEN_3031;
  wire  _GEN_3033 = 9'h1ff == out_iindex_1 ? _out_T_1122 : _GEN_3032;
  wire [31:0] _GEN_3035 = 9'h1 == out_iindex_1 ? 32'h380006f : 32'hc0006f;
  wire [31:0] _GEN_3036 = 9'h2 == out_iindex_1 ? 32'h440006f : _GEN_3035;
  wire [31:0] _GEN_3037 = 9'h3 == out_iindex_1 ? 32'hff0000f : _GEN_3036;
  wire [31:0] _GEN_3038 = 9'h4 == out_iindex_1 ? 32'h7b241073 : _GEN_3037;
  wire [31:0] _GEN_3039 = 9'h5 == out_iindex_1 ? 32'hf1402473 : _GEN_3038;
  wire [31:0] _GEN_3040 = 9'h6 == out_iindex_1 ? 32'h10802023 : _GEN_3039;
  wire [31:0] _GEN_3041 = 9'h7 == out_iindex_1 ? 32'h40044403 : _GEN_3040;
  wire [31:0] _GEN_3042 = 9'h8 == out_iindex_1 ? 32'h347413 : _GEN_3041;
  wire [31:0] _GEN_3043 = 9'h9 == out_iindex_1 ? 32'hfe0408e3 : _GEN_3042;
  wire [31:0] _GEN_3044 = 9'ha == out_iindex_1 ? 32'h147413 : _GEN_3043;
  wire [31:0] _GEN_3045 = 9'hb == out_iindex_1 ? 32'h40863 : _GEN_3044;
  wire [31:0] _GEN_3046 = 9'hc == out_iindex_1 ? 32'h7b202473 : _GEN_3045;
  wire [31:0] _GEN_3047 = 9'hd == out_iindex_1 ? 32'h10002223 : _GEN_3046;
  wire [31:0] _GEN_3048 = 9'he == out_iindex_1 ? 32'h30000067 : _GEN_3047;
  wire [31:0] _GEN_3049 = 9'hf == out_iindex_1 ? 32'hf1402473 : _GEN_3048;
  wire [31:0] _GEN_3050 = 9'h10 == out_iindex_1 ? 32'h10802423 : _GEN_3049;
  wire [31:0] _GEN_3051 = 9'h11 == out_iindex_1 ? 32'h7b202473 : _GEN_3050;
  wire [31:0] _GEN_3052 = 9'h12 == out_iindex_1 ? 32'h7b200073 : _GEN_3051;
  wire [31:0] _GEN_3053 = 9'h13 == out_iindex_1 ? 32'h10002623 : _GEN_3052;
  wire [31:0] _GEN_3054 = 9'h14 == out_iindex_1 ? 32'h100073 : _GEN_3053;
  wire [31:0] _GEN_3055 = 9'h15 == out_iindex_1 ? 32'h0 : _GEN_3054;
  wire [31:0] _GEN_3056 = 9'h16 == out_iindex_1 ? 32'h0 : _GEN_3055;
  wire [31:0] _GEN_3057 = 9'h17 == out_iindex_1 ? 32'h0 : _GEN_3056;
  wire [31:0] _GEN_3058 = 9'h18 == out_iindex_1 ? 32'h0 : _GEN_3057;
  wire [31:0] _GEN_3059 = 9'h19 == out_iindex_1 ? 32'h0 : _GEN_3058;
  wire [31:0] _GEN_3060 = 9'h1a == out_iindex_1 ? 32'h0 : _GEN_3059;
  wire [31:0] _GEN_3061 = 9'h1b == out_iindex_1 ? 32'h0 : _GEN_3060;
  wire [31:0] _GEN_3062 = 9'h1c == out_iindex_1 ? 32'h0 : _GEN_3061;
  wire [31:0] _GEN_3063 = 9'h1d == out_iindex_1 ? 32'h0 : _GEN_3062;
  wire [31:0] _GEN_3064 = 9'h1e == out_iindex_1 ? 32'h0 : _GEN_3063;
  wire [31:0] _GEN_3065 = 9'h1f == out_iindex_1 ? 32'h0 : _GEN_3064;
  wire [31:0] _GEN_3066 = 9'h20 == out_iindex_1 ? 32'h0 : _GEN_3065;
  wire [31:0] _GEN_3067 = 9'h21 == out_iindex_1 ? 32'h0 : _GEN_3066;
  wire [31:0] _GEN_3068 = 9'h22 == out_iindex_1 ? 32'h0 : _GEN_3067;
  wire [31:0] _GEN_3069 = 9'h23 == out_iindex_1 ? 32'h0 : _GEN_3068;
  wire [31:0] _GEN_3070 = 9'h24 == out_iindex_1 ? 32'h0 : _GEN_3069;
  wire [31:0] _GEN_3071 = 9'h25 == out_iindex_1 ? 32'h0 : _GEN_3070;
  wire [31:0] _GEN_3072 = 9'h26 == out_iindex_1 ? 32'h0 : _GEN_3071;
  wire [31:0] _GEN_3073 = 9'h27 == out_iindex_1 ? 32'h0 : _GEN_3072;
  wire [31:0] _GEN_3074 = 9'h28 == out_iindex_1 ? 32'h0 : _GEN_3073;
  wire [31:0] _GEN_3075 = 9'h29 == out_iindex_1 ? 32'h0 : _GEN_3074;
  wire [31:0] _GEN_3076 = 9'h2a == out_iindex_1 ? 32'h0 : _GEN_3075;
  wire [31:0] _GEN_3077 = 9'h2b == out_iindex_1 ? 32'h0 : _GEN_3076;
  wire [31:0] _GEN_3078 = 9'h2c == out_iindex_1 ? 32'h0 : _GEN_3077;
  wire [31:0] _GEN_3079 = 9'h2d == out_iindex_1 ? 32'h0 : _GEN_3078;
  wire [31:0] _GEN_3080 = 9'h2e == out_iindex_1 ? 32'h0 : _GEN_3079;
  wire [31:0] _GEN_3081 = 9'h2f == out_iindex_1 ? 32'h0 : _GEN_3080;
  wire [31:0] _GEN_3082 = 9'h30 == out_iindex_1 ? 32'h0 : _GEN_3081;
  wire [31:0] _GEN_3083 = 9'h31 == out_iindex_1 ? 32'h0 : _GEN_3082;
  wire [31:0] _GEN_3084 = 9'h32 == out_iindex_1 ? 32'h0 : _GEN_3083;
  wire [31:0] _GEN_3085 = 9'h33 == out_iindex_1 ? 32'h0 : _GEN_3084;
  wire [31:0] _GEN_3086 = 9'h34 == out_iindex_1 ? 32'h0 : _GEN_3085;
  wire [31:0] _GEN_3087 = 9'h35 == out_iindex_1 ? 32'h0 : _GEN_3086;
  wire [31:0] _GEN_3088 = 9'h36 == out_iindex_1 ? 32'h0 : _GEN_3087;
  wire [31:0] _GEN_3089 = 9'h37 == out_iindex_1 ? 32'h0 : _GEN_3088;
  wire [31:0] _GEN_3090 = 9'h38 == out_iindex_1 ? 32'h0 : _GEN_3089;
  wire [31:0] _GEN_3091 = 9'h39 == out_iindex_1 ? 32'h0 : _GEN_3090;
  wire [31:0] _GEN_3092 = 9'h3a == out_iindex_1 ? 32'h0 : _GEN_3091;
  wire [31:0] _GEN_3093 = 9'h3b == out_iindex_1 ? 32'h0 : _GEN_3092;
  wire [31:0] _GEN_3094 = 9'h3c == out_iindex_1 ? 32'h0 : _GEN_3093;
  wire [31:0] _GEN_3095 = 9'h3d == out_iindex_1 ? 32'h0 : _GEN_3094;
  wire [31:0] _GEN_3096 = 9'h3e == out_iindex_1 ? 32'h0 : _GEN_3095;
  wire [31:0] _GEN_3097 = 9'h3f == out_iindex_1 ? 32'h0 : _GEN_3096;
  wire [31:0] _GEN_3098 = 9'h40 == out_iindex_1 ? 32'h0 : _GEN_3097;
  wire [31:0] _GEN_3099 = 9'h41 == out_iindex_1 ? 32'h0 : _GEN_3098;
  wire [31:0] _GEN_3100 = 9'h42 == out_iindex_1 ? 32'h0 : _GEN_3099;
  wire [31:0] _GEN_3101 = 9'h43 == out_iindex_1 ? 32'h0 : _GEN_3100;
  wire [31:0] _GEN_3102 = 9'h44 == out_iindex_1 ? 32'h0 : _GEN_3101;
  wire [31:0] _GEN_3103 = 9'h45 == out_iindex_1 ? 32'h0 : _GEN_3102;
  wire [31:0] _GEN_3104 = 9'h46 == out_iindex_1 ? 32'h0 : _GEN_3103;
  wire [31:0] _GEN_3105 = 9'h47 == out_iindex_1 ? 32'h0 : _GEN_3104;
  wire [31:0] _GEN_3106 = 9'h48 == out_iindex_1 ? 32'h0 : _GEN_3105;
  wire [31:0] _GEN_3107 = 9'h49 == out_iindex_1 ? 32'h0 : _GEN_3106;
  wire [31:0] _GEN_3108 = 9'h4a == out_iindex_1 ? 32'h0 : _GEN_3107;
  wire [31:0] _GEN_3109 = 9'h4b == out_iindex_1 ? 32'h0 : _GEN_3108;
  wire [31:0] _GEN_3110 = 9'h4c == out_iindex_1 ? 32'h0 : _GEN_3109;
  wire [31:0] _GEN_3111 = 9'h4d == out_iindex_1 ? 32'h0 : _GEN_3110;
  wire [31:0] _GEN_3112 = 9'h4e == out_iindex_1 ? 32'h0 : _GEN_3111;
  wire [31:0] _GEN_3113 = 9'h4f == out_iindex_1 ? 32'h0 : _GEN_3112;
  wire [31:0] _GEN_3114 = 9'h50 == out_iindex_1 ? 32'h0 : _GEN_3113;
  wire [31:0] _GEN_3115 = 9'h51 == out_iindex_1 ? 32'h0 : _GEN_3114;
  wire [31:0] _GEN_3116 = 9'h52 == out_iindex_1 ? 32'h0 : _GEN_3115;
  wire [31:0] _GEN_3117 = 9'h53 == out_iindex_1 ? 32'h0 : _GEN_3116;
  wire [31:0] _GEN_3118 = 9'h54 == out_iindex_1 ? 32'h0 : _GEN_3117;
  wire [31:0] _GEN_3119 = 9'h55 == out_iindex_1 ? 32'h0 : _GEN_3118;
  wire [31:0] _GEN_3120 = 9'h56 == out_iindex_1 ? 32'h0 : _GEN_3119;
  wire [31:0] _GEN_3121 = 9'h57 == out_iindex_1 ? 32'h0 : _GEN_3120;
  wire [31:0] _GEN_3122 = 9'h58 == out_iindex_1 ? 32'h0 : _GEN_3121;
  wire [31:0] _GEN_3123 = 9'h59 == out_iindex_1 ? 32'h0 : _GEN_3122;
  wire [31:0] _GEN_3124 = 9'h5a == out_iindex_1 ? 32'h0 : _GEN_3123;
  wire [31:0] _GEN_3125 = 9'h5b == out_iindex_1 ? 32'h0 : _GEN_3124;
  wire [31:0] _GEN_3126 = 9'h5c == out_iindex_1 ? 32'h0 : _GEN_3125;
  wire [31:0] _GEN_3127 = 9'h5d == out_iindex_1 ? 32'h0 : _GEN_3126;
  wire [31:0] _GEN_3128 = 9'h5e == out_iindex_1 ? 32'h0 : _GEN_3127;
  wire [31:0] _GEN_3129 = 9'h5f == out_iindex_1 ? 32'h0 : _GEN_3128;
  wire [31:0] _GEN_3130 = 9'h60 == out_iindex_1 ? 32'h0 : _GEN_3129;
  wire [31:0] _GEN_3131 = 9'h61 == out_iindex_1 ? 32'h0 : _GEN_3130;
  wire [31:0] _GEN_3132 = 9'h62 == out_iindex_1 ? 32'h0 : _GEN_3131;
  wire [31:0] _GEN_3133 = 9'h63 == out_iindex_1 ? 32'h0 : _GEN_3132;
  wire [31:0] _GEN_3134 = 9'h64 == out_iindex_1 ? 32'h0 : _GEN_3133;
  wire [31:0] _GEN_3135 = 9'h65 == out_iindex_1 ? 32'h0 : _GEN_3134;
  wire [31:0] _GEN_3136 = 9'h66 == out_iindex_1 ? 32'h0 : _GEN_3135;
  wire [31:0] _GEN_3137 = 9'h67 == out_iindex_1 ? 32'h0 : _GEN_3136;
  wire [31:0] _GEN_3138 = 9'h68 == out_iindex_1 ? 32'h0 : _GEN_3137;
  wire [31:0] _GEN_3139 = 9'h69 == out_iindex_1 ? 32'h0 : _GEN_3138;
  wire [31:0] _GEN_3140 = 9'h6a == out_iindex_1 ? 32'h0 : _GEN_3139;
  wire [31:0] _GEN_3141 = 9'h6b == out_iindex_1 ? 32'h0 : _GEN_3140;
  wire [31:0] _GEN_3142 = 9'h6c == out_iindex_1 ? 32'h0 : _GEN_3141;
  wire [31:0] _GEN_3143 = 9'h6d == out_iindex_1 ? 32'h0 : _GEN_3142;
  wire [31:0] _GEN_3144 = 9'h6e == out_iindex_1 ? 32'h0 : _GEN_3143;
  wire [31:0] _GEN_3145 = 9'h6f == out_iindex_1 ? 32'h0 : _GEN_3144;
  wire [31:0] _GEN_3146 = 9'h70 == out_iindex_1 ? 32'h0 : _GEN_3145;
  wire [31:0] _GEN_3147 = 9'h71 == out_iindex_1 ? 32'h0 : _GEN_3146;
  wire [31:0] _GEN_3148 = 9'h72 == out_iindex_1 ? 32'h0 : _GEN_3147;
  wire [31:0] _GEN_3149 = 9'h73 == out_iindex_1 ? 32'h0 : _GEN_3148;
  wire [31:0] _GEN_3150 = 9'h74 == out_iindex_1 ? 32'h0 : _GEN_3149;
  wire [31:0] _GEN_3151 = 9'h75 == out_iindex_1 ? 32'h0 : _GEN_3150;
  wire [31:0] _GEN_3152 = 9'h76 == out_iindex_1 ? 32'h0 : _GEN_3151;
  wire [31:0] _GEN_3153 = 9'h77 == out_iindex_1 ? 32'h0 : _GEN_3152;
  wire [31:0] _GEN_3154 = 9'h78 == out_iindex_1 ? 32'h0 : _GEN_3153;
  wire [31:0] _GEN_3155 = 9'h79 == out_iindex_1 ? 32'h0 : _GEN_3154;
  wire [31:0] _GEN_3156 = 9'h7a == out_iindex_1 ? 32'h0 : _GEN_3155;
  wire [31:0] _GEN_3157 = 9'h7b == out_iindex_1 ? 32'h0 : _GEN_3156;
  wire [31:0] _GEN_3158 = 9'h7c == out_iindex_1 ? 32'h0 : _GEN_3157;
  wire [31:0] _GEN_3159 = 9'h7d == out_iindex_1 ? 32'h0 : _GEN_3158;
  wire [31:0] _GEN_3160 = 9'h7e == out_iindex_1 ? 32'h0 : _GEN_3159;
  wire [31:0] _GEN_3161 = 9'h7f == out_iindex_1 ? 32'h0 : _GEN_3160;
  wire [31:0] _GEN_3162 = 9'h80 == out_iindex_1 ? 32'h0 : _GEN_3161;
  wire [31:0] _GEN_3163 = 9'h81 == out_iindex_1 ? 32'h0 : _GEN_3162;
  wire [31:0] _GEN_3164 = 9'h82 == out_iindex_1 ? 32'h0 : _GEN_3163;
  wire [31:0] _GEN_3165 = 9'h83 == out_iindex_1 ? 32'h0 : _GEN_3164;
  wire [31:0] _GEN_3166 = 9'h84 == out_iindex_1 ? 32'h0 : _GEN_3165;
  wire [31:0] _GEN_3167 = 9'h85 == out_iindex_1 ? 32'h0 : _GEN_3166;
  wire [31:0] _GEN_3168 = 9'h86 == out_iindex_1 ? 32'h0 : _GEN_3167;
  wire [31:0] _GEN_3169 = 9'h87 == out_iindex_1 ? 32'h0 : _GEN_3168;
  wire [31:0] _GEN_3170 = 9'h88 == out_iindex_1 ? 32'h0 : _GEN_3169;
  wire [31:0] _GEN_3171 = 9'h89 == out_iindex_1 ? 32'h0 : _GEN_3170;
  wire [31:0] _GEN_3172 = 9'h8a == out_iindex_1 ? 32'h0 : _GEN_3171;
  wire [31:0] _GEN_3173 = 9'h8b == out_iindex_1 ? 32'h0 : _GEN_3172;
  wire [31:0] _GEN_3174 = 9'h8c == out_iindex_1 ? 32'h0 : _GEN_3173;
  wire [31:0] _GEN_3175 = 9'h8d == out_iindex_1 ? 32'h0 : _GEN_3174;
  wire [31:0] _GEN_3176 = 9'h8e == out_iindex_1 ? 32'h0 : _GEN_3175;
  wire [31:0] _GEN_3177 = 9'h8f == out_iindex_1 ? 32'h0 : _GEN_3176;
  wire [31:0] _GEN_3178 = 9'h90 == out_iindex_1 ? 32'h0 : _GEN_3177;
  wire [31:0] _GEN_3179 = 9'h91 == out_iindex_1 ? 32'h0 : _GEN_3178;
  wire [31:0] _GEN_3180 = 9'h92 == out_iindex_1 ? 32'h0 : _GEN_3179;
  wire [31:0] _GEN_3181 = 9'h93 == out_iindex_1 ? 32'h0 : _GEN_3180;
  wire [31:0] _GEN_3182 = 9'h94 == out_iindex_1 ? 32'h0 : _GEN_3181;
  wire [31:0] _GEN_3183 = 9'h95 == out_iindex_1 ? 32'h0 : _GEN_3182;
  wire [31:0] _GEN_3184 = 9'h96 == out_iindex_1 ? 32'h0 : _GEN_3183;
  wire [31:0] _GEN_3185 = 9'h97 == out_iindex_1 ? 32'h0 : _GEN_3184;
  wire [31:0] _GEN_3186 = 9'h98 == out_iindex_1 ? 32'h0 : _GEN_3185;
  wire [31:0] _GEN_3187 = 9'h99 == out_iindex_1 ? 32'h0 : _GEN_3186;
  wire [31:0] _GEN_3188 = 9'h9a == out_iindex_1 ? 32'h0 : _GEN_3187;
  wire [31:0] _GEN_3189 = 9'h9b == out_iindex_1 ? 32'h0 : _GEN_3188;
  wire [31:0] _GEN_3190 = 9'h9c == out_iindex_1 ? 32'h0 : _GEN_3189;
  wire [31:0] _GEN_3191 = 9'h9d == out_iindex_1 ? 32'h0 : _GEN_3190;
  wire [31:0] _GEN_3192 = 9'h9e == out_iindex_1 ? 32'h0 : _GEN_3191;
  wire [31:0] _GEN_3193 = 9'h9f == out_iindex_1 ? 32'h0 : _GEN_3192;
  wire [31:0] _GEN_3194 = 9'ha0 == out_iindex_1 ? 32'h0 : _GEN_3193;
  wire [31:0] _GEN_3195 = 9'ha1 == out_iindex_1 ? 32'h0 : _GEN_3194;
  wire [31:0] _GEN_3196 = 9'ha2 == out_iindex_1 ? 32'h0 : _GEN_3195;
  wire [31:0] _GEN_3197 = 9'ha3 == out_iindex_1 ? 32'h0 : _GEN_3196;
  wire [31:0] _GEN_3198 = 9'ha4 == out_iindex_1 ? 32'h0 : _GEN_3197;
  wire [31:0] _GEN_3199 = 9'ha5 == out_iindex_1 ? 32'h0 : _GEN_3198;
  wire [31:0] _GEN_3200 = 9'ha6 == out_iindex_1 ? 32'h0 : _GEN_3199;
  wire [31:0] _GEN_3201 = 9'ha7 == out_iindex_1 ? 32'h0 : _GEN_3200;
  wire [31:0] _GEN_3202 = 9'ha8 == out_iindex_1 ? 32'h0 : _GEN_3201;
  wire [31:0] _GEN_3203 = 9'ha9 == out_iindex_1 ? 32'h0 : _GEN_3202;
  wire [31:0] _GEN_3204 = 9'haa == out_iindex_1 ? 32'h0 : _GEN_3203;
  wire [31:0] _GEN_3205 = 9'hab == out_iindex_1 ? 32'h0 : _GEN_3204;
  wire [31:0] _GEN_3206 = 9'hac == out_iindex_1 ? 32'h0 : _GEN_3205;
  wire [31:0] _GEN_3207 = 9'had == out_iindex_1 ? 32'h0 : _GEN_3206;
  wire [31:0] _GEN_3208 = 9'hae == out_iindex_1 ? 32'h0 : _GEN_3207;
  wire [31:0] _GEN_3209 = 9'haf == out_iindex_1 ? 32'h0 : _GEN_3208;
  wire [31:0] _GEN_3210 = 9'hb0 == out_iindex_1 ? 32'h0 : _GEN_3209;
  wire [31:0] _GEN_3211 = 9'hb1 == out_iindex_1 ? 32'h0 : _GEN_3210;
  wire [31:0] _GEN_3212 = 9'hb2 == out_iindex_1 ? 32'h0 : _GEN_3211;
  wire [31:0] _GEN_3213 = 9'hb3 == out_iindex_1 ? 32'h0 : _GEN_3212;
  wire [31:0] _GEN_3214 = 9'hb4 == out_iindex_1 ? 32'h0 : _GEN_3213;
  wire [31:0] _GEN_3215 = 9'hb5 == out_iindex_1 ? 32'h0 : _GEN_3214;
  wire [31:0] _GEN_3216 = 9'hb6 == out_iindex_1 ? 32'h0 : _GEN_3215;
  wire [31:0] _GEN_3217 = 9'hb7 == out_iindex_1 ? 32'h0 : _GEN_3216;
  wire [31:0] _GEN_3218 = 9'hb8 == out_iindex_1 ? 32'h0 : _GEN_3217;
  wire [31:0] _GEN_3219 = 9'hb9 == out_iindex_1 ? 32'h0 : _GEN_3218;
  wire [31:0] _GEN_3220 = 9'hba == out_iindex_1 ? 32'h0 : _GEN_3219;
  wire [31:0] _GEN_3221 = 9'hbb == out_iindex_1 ? 32'h0 : _GEN_3220;
  wire [31:0] _GEN_3222 = 9'hbc == out_iindex_1 ? 32'h0 : _GEN_3221;
  wire [31:0] _GEN_3223 = 9'hbd == out_iindex_1 ? 32'h0 : _GEN_3222;
  wire [31:0] _GEN_3224 = 9'hbe == out_iindex_1 ? 32'h0 : _GEN_3223;
  wire [31:0] _GEN_3225 = 9'hbf == out_iindex_1 ? 32'h0 : _GEN_3224;
  wire [31:0] _GEN_3226 = 9'hc0 == out_iindex_1 ? 32'h380006f : _GEN_3225;
  wire [31:0] _GEN_3227 = 9'hc1 == out_iindex_1 ? 32'h0 : _GEN_3226;
  wire [31:0] _GEN_3228 = 9'hc2 == out_iindex_1 ? 32'h0 : _GEN_3227;
  wire [31:0] _GEN_3229 = 9'hc3 == out_iindex_1 ? 32'h0 : _GEN_3228;
  wire [31:0] _GEN_3230 = 9'hc4 == out_iindex_1 ? 32'h0 : _GEN_3229;
  wire [31:0] _GEN_3231 = 9'hc5 == out_iindex_1 ? 32'h0 : _GEN_3230;
  wire [31:0] _GEN_3232 = 9'hc6 == out_iindex_1 ? 32'h0 : _GEN_3231;
  wire [31:0] _GEN_3233 = 9'hc7 == out_iindex_1 ? 32'h0 : _GEN_3232;
  wire [31:0] _GEN_3234 = 9'hc8 == out_iindex_1 ? 32'h0 : _GEN_3233;
  wire [31:0] _GEN_3235 = 9'hc9 == out_iindex_1 ? 32'h0 : _GEN_3234;
  wire [31:0] _GEN_3236 = 9'hca == out_iindex_1 ? 32'h0 : _GEN_3235;
  wire [31:0] _GEN_3237 = 9'hcb == out_iindex_1 ? 32'h0 : _GEN_3236;
  wire [31:0] _GEN_3238 = 9'hcc == out_iindex_1 ? 32'h0 : _GEN_3237;
  wire [31:0] _GEN_3239 = 9'hcd == out_iindex_1 ? 32'h0 : _GEN_3238;
  wire [31:0] _GEN_3240 = 9'hce == out_iindex_1 ? abstractGeneratedMem_0 : _GEN_3239;
  wire [31:0] _GEN_3241 = 9'hcf == out_iindex_1 ? abstractGeneratedMem_1 : _GEN_3240;
  wire [31:0] _GEN_3242 = 9'hd0 == out_iindex_1 ? out_prepend_22 : _GEN_3241;
  wire [31:0] _GEN_3243 = 9'hd1 == out_iindex_1 ? out_prepend_16 : _GEN_3242;
  wire [31:0] _GEN_3244 = 9'hd2 == out_iindex_1 ? out_prepend_25 : _GEN_3243;
  wire [31:0] _GEN_3245 = 9'hd3 == out_iindex_1 ? out_prepend_61 : _GEN_3244;
  wire [31:0] _GEN_3246 = 9'hd4 == out_iindex_1 ? out_prepend_70 : _GEN_3245;
  wire [31:0] _GEN_3247 = 9'hd5 == out_iindex_1 ? out_prepend_7 : _GEN_3246;
  wire [31:0] _GEN_3248 = 9'hd6 == out_iindex_1 ? out_prepend_13 : _GEN_3247;
  wire [31:0] _GEN_3249 = 9'hd7 == out_iindex_1 ? out_prepend_58 : _GEN_3248;
  wire [31:0] _GEN_3250 = 9'hd8 == out_iindex_1 ? out_prepend_67 : _GEN_3249;
  wire [31:0] _GEN_3251 = 9'hd9 == out_iindex_1 ? out_prepend_19 : _GEN_3250;
  wire [31:0] _GEN_3252 = 9'hda == out_iindex_1 ? out_prepend_2 : _GEN_3251;
  wire [31:0] _GEN_3253 = 9'hdb == out_iindex_1 ? out_prepend_64 : _GEN_3252;
  wire [31:0] _GEN_3254 = 9'hdc == out_iindex_1 ? out_prepend_55 : _GEN_3253;
  wire [31:0] _GEN_3255 = 9'hdd == out_iindex_1 ? out_prepend_28 : _GEN_3254;
  wire [31:0] _GEN_3256 = 9'hde == out_iindex_1 ? out_prepend_10 : _GEN_3255;
  wire [31:0] _GEN_3257 = 9'hdf == out_iindex_1 ? out_prepend_76 : _GEN_3256;
  wire [31:0] _GEN_3258 = 9'he0 == out_iindex_1 ? out_prepend_73 : _GEN_3257;
  wire [31:0] _GEN_3259 = 9'he1 == out_iindex_1 ? 32'h0 : _GEN_3258;
  wire [31:0] _GEN_3260 = 9'he2 == out_iindex_1 ? 32'h0 : _GEN_3259;
  wire [31:0] _GEN_3261 = 9'he3 == out_iindex_1 ? 32'h0 : _GEN_3260;
  wire [31:0] _GEN_3262 = 9'he4 == out_iindex_1 ? 32'h0 : _GEN_3261;
  wire [31:0] _GEN_3263 = 9'he5 == out_iindex_1 ? 32'h0 : _GEN_3262;
  wire [31:0] _GEN_3264 = 9'he6 == out_iindex_1 ? 32'h0 : _GEN_3263;
  wire [31:0] _GEN_3265 = 9'he7 == out_iindex_1 ? 32'h0 : _GEN_3264;
  wire [31:0] _GEN_3266 = 9'he8 == out_iindex_1 ? 32'h0 : _GEN_3265;
  wire [31:0] _GEN_3267 = 9'he9 == out_iindex_1 ? 32'h0 : _GEN_3266;
  wire [31:0] _GEN_3268 = 9'hea == out_iindex_1 ? 32'h0 : _GEN_3267;
  wire [31:0] _GEN_3269 = 9'heb == out_iindex_1 ? 32'h0 : _GEN_3268;
  wire [31:0] _GEN_3270 = 9'hec == out_iindex_1 ? 32'h0 : _GEN_3269;
  wire [31:0] _GEN_3271 = 9'hed == out_iindex_1 ? 32'h0 : _GEN_3270;
  wire [31:0] _GEN_3272 = 9'hee == out_iindex_1 ? 32'h0 : _GEN_3271;
  wire [31:0] _GEN_3273 = 9'hef == out_iindex_1 ? 32'h0 : _GEN_3272;
  wire [31:0] _GEN_3274 = 9'hf0 == out_iindex_1 ? 32'h0 : _GEN_3273;
  wire [31:0] _GEN_3275 = 9'hf1 == out_iindex_1 ? 32'h0 : _GEN_3274;
  wire [31:0] _GEN_3276 = 9'hf2 == out_iindex_1 ? 32'h0 : _GEN_3275;
  wire [31:0] _GEN_3277 = 9'hf3 == out_iindex_1 ? 32'h0 : _GEN_3276;
  wire [31:0] _GEN_3278 = 9'hf4 == out_iindex_1 ? 32'h0 : _GEN_3277;
  wire [31:0] _GEN_3279 = 9'hf5 == out_iindex_1 ? 32'h0 : _GEN_3278;
  wire [31:0] _GEN_3280 = 9'hf6 == out_iindex_1 ? 32'h0 : _GEN_3279;
  wire [31:0] _GEN_3281 = 9'hf7 == out_iindex_1 ? 32'h0 : _GEN_3280;
  wire [31:0] _GEN_3282 = 9'hf8 == out_iindex_1 ? 32'h0 : _GEN_3281;
  wire [31:0] _GEN_3283 = 9'hf9 == out_iindex_1 ? 32'h0 : _GEN_3282;
  wire [31:0] _GEN_3284 = 9'hfa == out_iindex_1 ? 32'h0 : _GEN_3283;
  wire [31:0] _GEN_3285 = 9'hfb == out_iindex_1 ? 32'h0 : _GEN_3284;
  wire [31:0] _GEN_3286 = 9'hfc == out_iindex_1 ? 32'h0 : _GEN_3285;
  wire [31:0] _GEN_3287 = 9'hfd == out_iindex_1 ? 32'h0 : _GEN_3286;
  wire [31:0] _GEN_3288 = 9'hfe == out_iindex_1 ? 32'h0 : _GEN_3287;
  wire [31:0] _GEN_3289 = 9'hff == out_iindex_1 ? 32'h0 : _GEN_3288;
  wire [31:0] _GEN_3290 = 9'h100 == out_iindex_1 ? out_prepend_79 : _GEN_3289;
  wire [31:0] _GEN_3291 = 9'h101 == out_iindex_1 ? out_prepend_79 : _GEN_3290;
  wire [31:0] _GEN_3292 = 9'h102 == out_iindex_1 ? out_prepend_79 : _GEN_3291;
  wire [31:0] _GEN_3293 = 9'h103 == out_iindex_1 ? out_prepend_79 : _GEN_3292;
  wire [31:0] _GEN_3294 = 9'h104 == out_iindex_1 ? out_prepend_79 : _GEN_3293;
  wire [31:0] _GEN_3295 = 9'h105 == out_iindex_1 ? out_prepend_79 : _GEN_3294;
  wire [31:0] _GEN_3296 = 9'h106 == out_iindex_1 ? out_prepend_79 : _GEN_3295;
  wire [31:0] _GEN_3297 = 9'h107 == out_iindex_1 ? out_prepend_79 : _GEN_3296;
  wire [31:0] _GEN_3298 = 9'h108 == out_iindex_1 ? out_prepend_79 : _GEN_3297;
  wire [31:0] _GEN_3299 = 9'h109 == out_iindex_1 ? out_prepend_79 : _GEN_3298;
  wire [31:0] _GEN_3300 = 9'h10a == out_iindex_1 ? out_prepend_79 : _GEN_3299;
  wire [31:0] _GEN_3301 = 9'h10b == out_iindex_1 ? out_prepend_79 : _GEN_3300;
  wire [31:0] _GEN_3302 = 9'h10c == out_iindex_1 ? out_prepend_79 : _GEN_3301;
  wire [31:0] _GEN_3303 = 9'h10d == out_iindex_1 ? out_prepend_79 : _GEN_3302;
  wire [31:0] _GEN_3304 = 9'h10e == out_iindex_1 ? out_prepend_79 : _GEN_3303;
  wire [31:0] _GEN_3305 = 9'h10f == out_iindex_1 ? out_prepend_79 : _GEN_3304;
  wire [31:0] _GEN_3306 = 9'h110 == out_iindex_1 ? out_prepend_79 : _GEN_3305;
  wire [31:0] _GEN_3307 = 9'h111 == out_iindex_1 ? out_prepend_79 : _GEN_3306;
  wire [31:0] _GEN_3308 = 9'h112 == out_iindex_1 ? out_prepend_79 : _GEN_3307;
  wire [31:0] _GEN_3309 = 9'h113 == out_iindex_1 ? out_prepend_79 : _GEN_3308;
  wire [31:0] _GEN_3310 = 9'h114 == out_iindex_1 ? out_prepend_79 : _GEN_3309;
  wire [31:0] _GEN_3311 = 9'h115 == out_iindex_1 ? out_prepend_79 : _GEN_3310;
  wire [31:0] _GEN_3312 = 9'h116 == out_iindex_1 ? out_prepend_79 : _GEN_3311;
  wire [31:0] _GEN_3313 = 9'h117 == out_iindex_1 ? out_prepend_79 : _GEN_3312;
  wire [31:0] _GEN_3314 = 9'h118 == out_iindex_1 ? out_prepend_79 : _GEN_3313;
  wire [31:0] _GEN_3315 = 9'h119 == out_iindex_1 ? out_prepend_79 : _GEN_3314;
  wire [31:0] _GEN_3316 = 9'h11a == out_iindex_1 ? out_prepend_79 : _GEN_3315;
  wire [31:0] _GEN_3317 = 9'h11b == out_iindex_1 ? out_prepend_79 : _GEN_3316;
  wire [31:0] _GEN_3318 = 9'h11c == out_iindex_1 ? out_prepend_79 : _GEN_3317;
  wire [31:0] _GEN_3319 = 9'h11d == out_iindex_1 ? out_prepend_79 : _GEN_3318;
  wire [31:0] _GEN_3320 = 9'h11e == out_iindex_1 ? out_prepend_79 : _GEN_3319;
  wire [31:0] _GEN_3321 = 9'h11f == out_iindex_1 ? out_prepend_79 : _GEN_3320;
  wire [31:0] _GEN_3322 = 9'h120 == out_iindex_1 ? out_prepend_79 : _GEN_3321;
  wire [31:0] _GEN_3323 = 9'h121 == out_iindex_1 ? out_prepend_79 : _GEN_3322;
  wire [31:0] _GEN_3324 = 9'h122 == out_iindex_1 ? out_prepend_79 : _GEN_3323;
  wire [31:0] _GEN_3325 = 9'h123 == out_iindex_1 ? out_prepend_79 : _GEN_3324;
  wire [31:0] _GEN_3326 = 9'h124 == out_iindex_1 ? out_prepend_79 : _GEN_3325;
  wire [31:0] _GEN_3327 = 9'h125 == out_iindex_1 ? out_prepend_79 : _GEN_3326;
  wire [31:0] _GEN_3328 = 9'h126 == out_iindex_1 ? out_prepend_79 : _GEN_3327;
  wire [31:0] _GEN_3329 = 9'h127 == out_iindex_1 ? out_prepend_79 : _GEN_3328;
  wire [31:0] _GEN_3330 = 9'h128 == out_iindex_1 ? out_prepend_79 : _GEN_3329;
  wire [31:0] _GEN_3331 = 9'h129 == out_iindex_1 ? out_prepend_79 : _GEN_3330;
  wire [31:0] _GEN_3332 = 9'h12a == out_iindex_1 ? out_prepend_79 : _GEN_3331;
  wire [31:0] _GEN_3333 = 9'h12b == out_iindex_1 ? out_prepend_79 : _GEN_3332;
  wire [31:0] _GEN_3334 = 9'h12c == out_iindex_1 ? out_prepend_79 : _GEN_3333;
  wire [31:0] _GEN_3335 = 9'h12d == out_iindex_1 ? out_prepend_79 : _GEN_3334;
  wire [31:0] _GEN_3336 = 9'h12e == out_iindex_1 ? out_prepend_79 : _GEN_3335;
  wire [31:0] _GEN_3337 = 9'h12f == out_iindex_1 ? out_prepend_79 : _GEN_3336;
  wire [31:0] _GEN_3338 = 9'h130 == out_iindex_1 ? out_prepend_79 : _GEN_3337;
  wire [31:0] _GEN_3339 = 9'h131 == out_iindex_1 ? out_prepend_79 : _GEN_3338;
  wire [31:0] _GEN_3340 = 9'h132 == out_iindex_1 ? out_prepend_79 : _GEN_3339;
  wire [31:0] _GEN_3341 = 9'h133 == out_iindex_1 ? out_prepend_79 : _GEN_3340;
  wire [31:0] _GEN_3342 = 9'h134 == out_iindex_1 ? out_prepend_79 : _GEN_3341;
  wire [31:0] _GEN_3343 = 9'h135 == out_iindex_1 ? out_prepend_79 : _GEN_3342;
  wire [31:0] _GEN_3344 = 9'h136 == out_iindex_1 ? out_prepend_79 : _GEN_3343;
  wire [31:0] _GEN_3345 = 9'h137 == out_iindex_1 ? out_prepend_79 : _GEN_3344;
  wire [31:0] _GEN_3346 = 9'h138 == out_iindex_1 ? out_prepend_79 : _GEN_3345;
  wire [31:0] _GEN_3347 = 9'h139 == out_iindex_1 ? out_prepend_79 : _GEN_3346;
  wire [31:0] _GEN_3348 = 9'h13a == out_iindex_1 ? out_prepend_79 : _GEN_3347;
  wire [31:0] _GEN_3349 = 9'h13b == out_iindex_1 ? out_prepend_79 : _GEN_3348;
  wire [31:0] _GEN_3350 = 9'h13c == out_iindex_1 ? out_prepend_79 : _GEN_3349;
  wire [31:0] _GEN_3351 = 9'h13d == out_iindex_1 ? out_prepend_79 : _GEN_3350;
  wire [31:0] _GEN_3352 = 9'h13e == out_iindex_1 ? out_prepend_79 : _GEN_3351;
  wire [31:0] _GEN_3353 = 9'h13f == out_iindex_1 ? out_prepend_79 : _GEN_3352;
  wire [31:0] _GEN_3354 = 9'h140 == out_iindex_1 ? out_prepend_79 : _GEN_3353;
  wire [31:0] _GEN_3355 = 9'h141 == out_iindex_1 ? out_prepend_79 : _GEN_3354;
  wire [31:0] _GEN_3356 = 9'h142 == out_iindex_1 ? out_prepend_79 : _GEN_3355;
  wire [31:0] _GEN_3357 = 9'h143 == out_iindex_1 ? out_prepend_79 : _GEN_3356;
  wire [31:0] _GEN_3358 = 9'h144 == out_iindex_1 ? out_prepend_79 : _GEN_3357;
  wire [31:0] _GEN_3359 = 9'h145 == out_iindex_1 ? out_prepend_79 : _GEN_3358;
  wire [31:0] _GEN_3360 = 9'h146 == out_iindex_1 ? out_prepend_79 : _GEN_3359;
  wire [31:0] _GEN_3361 = 9'h147 == out_iindex_1 ? out_prepend_79 : _GEN_3360;
  wire [31:0] _GEN_3362 = 9'h148 == out_iindex_1 ? out_prepend_79 : _GEN_3361;
  wire [31:0] _GEN_3363 = 9'h149 == out_iindex_1 ? out_prepend_79 : _GEN_3362;
  wire [31:0] _GEN_3364 = 9'h14a == out_iindex_1 ? out_prepend_79 : _GEN_3363;
  wire [31:0] _GEN_3365 = 9'h14b == out_iindex_1 ? out_prepend_79 : _GEN_3364;
  wire [31:0] _GEN_3366 = 9'h14c == out_iindex_1 ? out_prepend_79 : _GEN_3365;
  wire [31:0] _GEN_3367 = 9'h14d == out_iindex_1 ? out_prepend_79 : _GEN_3366;
  wire [31:0] _GEN_3368 = 9'h14e == out_iindex_1 ? out_prepend_79 : _GEN_3367;
  wire [31:0] _GEN_3369 = 9'h14f == out_iindex_1 ? out_prepend_79 : _GEN_3368;
  wire [31:0] _GEN_3370 = 9'h150 == out_iindex_1 ? out_prepend_79 : _GEN_3369;
  wire [31:0] _GEN_3371 = 9'h151 == out_iindex_1 ? out_prepend_79 : _GEN_3370;
  wire [31:0] _GEN_3372 = 9'h152 == out_iindex_1 ? out_prepend_79 : _GEN_3371;
  wire [31:0] _GEN_3373 = 9'h153 == out_iindex_1 ? out_prepend_79 : _GEN_3372;
  wire [31:0] _GEN_3374 = 9'h154 == out_iindex_1 ? out_prepend_79 : _GEN_3373;
  wire [31:0] _GEN_3375 = 9'h155 == out_iindex_1 ? out_prepend_79 : _GEN_3374;
  wire [31:0] _GEN_3376 = 9'h156 == out_iindex_1 ? out_prepend_79 : _GEN_3375;
  wire [31:0] _GEN_3377 = 9'h157 == out_iindex_1 ? out_prepend_79 : _GEN_3376;
  wire [31:0] _GEN_3378 = 9'h158 == out_iindex_1 ? out_prepend_79 : _GEN_3377;
  wire [31:0] _GEN_3379 = 9'h159 == out_iindex_1 ? out_prepend_79 : _GEN_3378;
  wire [31:0] _GEN_3380 = 9'h15a == out_iindex_1 ? out_prepend_79 : _GEN_3379;
  wire [31:0] _GEN_3381 = 9'h15b == out_iindex_1 ? out_prepend_79 : _GEN_3380;
  wire [31:0] _GEN_3382 = 9'h15c == out_iindex_1 ? out_prepend_79 : _GEN_3381;
  wire [31:0] _GEN_3383 = 9'h15d == out_iindex_1 ? out_prepend_79 : _GEN_3382;
  wire [31:0] _GEN_3384 = 9'h15e == out_iindex_1 ? out_prepend_79 : _GEN_3383;
  wire [31:0] _GEN_3385 = 9'h15f == out_iindex_1 ? out_prepend_79 : _GEN_3384;
  wire [31:0] _GEN_3386 = 9'h160 == out_iindex_1 ? out_prepend_79 : _GEN_3385;
  wire [31:0] _GEN_3387 = 9'h161 == out_iindex_1 ? out_prepend_79 : _GEN_3386;
  wire [31:0] _GEN_3388 = 9'h162 == out_iindex_1 ? out_prepend_79 : _GEN_3387;
  wire [31:0] _GEN_3389 = 9'h163 == out_iindex_1 ? out_prepend_79 : _GEN_3388;
  wire [31:0] _GEN_3390 = 9'h164 == out_iindex_1 ? out_prepend_79 : _GEN_3389;
  wire [31:0] _GEN_3391 = 9'h165 == out_iindex_1 ? out_prepend_79 : _GEN_3390;
  wire [31:0] _GEN_3392 = 9'h166 == out_iindex_1 ? out_prepend_79 : _GEN_3391;
  wire [31:0] _GEN_3393 = 9'h167 == out_iindex_1 ? out_prepend_79 : _GEN_3392;
  wire [31:0] _GEN_3394 = 9'h168 == out_iindex_1 ? out_prepend_79 : _GEN_3393;
  wire [31:0] _GEN_3395 = 9'h169 == out_iindex_1 ? out_prepend_79 : _GEN_3394;
  wire [31:0] _GEN_3396 = 9'h16a == out_iindex_1 ? out_prepend_79 : _GEN_3395;
  wire [31:0] _GEN_3397 = 9'h16b == out_iindex_1 ? out_prepend_79 : _GEN_3396;
  wire [31:0] _GEN_3398 = 9'h16c == out_iindex_1 ? out_prepend_79 : _GEN_3397;
  wire [31:0] _GEN_3399 = 9'h16d == out_iindex_1 ? out_prepend_79 : _GEN_3398;
  wire [31:0] _GEN_3400 = 9'h16e == out_iindex_1 ? out_prepend_79 : _GEN_3399;
  wire [31:0] _GEN_3401 = 9'h16f == out_iindex_1 ? out_prepend_79 : _GEN_3400;
  wire [31:0] _GEN_3402 = 9'h170 == out_iindex_1 ? out_prepend_79 : _GEN_3401;
  wire [31:0] _GEN_3403 = 9'h171 == out_iindex_1 ? out_prepend_79 : _GEN_3402;
  wire [31:0] _GEN_3404 = 9'h172 == out_iindex_1 ? out_prepend_79 : _GEN_3403;
  wire [31:0] _GEN_3405 = 9'h173 == out_iindex_1 ? out_prepend_79 : _GEN_3404;
  wire [31:0] _GEN_3406 = 9'h174 == out_iindex_1 ? out_prepend_79 : _GEN_3405;
  wire [31:0] _GEN_3407 = 9'h175 == out_iindex_1 ? out_prepend_79 : _GEN_3406;
  wire [31:0] _GEN_3408 = 9'h176 == out_iindex_1 ? out_prepend_79 : _GEN_3407;
  wire [31:0] _GEN_3409 = 9'h177 == out_iindex_1 ? out_prepend_79 : _GEN_3408;
  wire [31:0] _GEN_3410 = 9'h178 == out_iindex_1 ? out_prepend_79 : _GEN_3409;
  wire [31:0] _GEN_3411 = 9'h179 == out_iindex_1 ? out_prepend_79 : _GEN_3410;
  wire [31:0] _GEN_3412 = 9'h17a == out_iindex_1 ? out_prepend_79 : _GEN_3411;
  wire [31:0] _GEN_3413 = 9'h17b == out_iindex_1 ? out_prepend_79 : _GEN_3412;
  wire [31:0] _GEN_3414 = 9'h17c == out_iindex_1 ? out_prepend_79 : _GEN_3413;
  wire [31:0] _GEN_3415 = 9'h17d == out_iindex_1 ? out_prepend_79 : _GEN_3414;
  wire [31:0] _GEN_3416 = 9'h17e == out_iindex_1 ? out_prepend_79 : _GEN_3415;
  wire [31:0] _GEN_3417 = 9'h17f == out_iindex_1 ? out_prepend_79 : _GEN_3416;
  wire [31:0] _GEN_3418 = 9'h180 == out_iindex_1 ? out_prepend_79 : _GEN_3417;
  wire [31:0] _GEN_3419 = 9'h181 == out_iindex_1 ? out_prepend_79 : _GEN_3418;
  wire [31:0] _GEN_3420 = 9'h182 == out_iindex_1 ? out_prepend_79 : _GEN_3419;
  wire [31:0] _GEN_3421 = 9'h183 == out_iindex_1 ? out_prepend_79 : _GEN_3420;
  wire [31:0] _GEN_3422 = 9'h184 == out_iindex_1 ? out_prepend_79 : _GEN_3421;
  wire [31:0] _GEN_3423 = 9'h185 == out_iindex_1 ? out_prepend_79 : _GEN_3422;
  wire [31:0] _GEN_3424 = 9'h186 == out_iindex_1 ? out_prepend_79 : _GEN_3423;
  wire [31:0] _GEN_3425 = 9'h187 == out_iindex_1 ? out_prepend_79 : _GEN_3424;
  wire [31:0] _GEN_3426 = 9'h188 == out_iindex_1 ? out_prepend_79 : _GEN_3425;
  wire [31:0] _GEN_3427 = 9'h189 == out_iindex_1 ? out_prepend_79 : _GEN_3426;
  wire [31:0] _GEN_3428 = 9'h18a == out_iindex_1 ? out_prepend_79 : _GEN_3427;
  wire [31:0] _GEN_3429 = 9'h18b == out_iindex_1 ? out_prepend_79 : _GEN_3428;
  wire [31:0] _GEN_3430 = 9'h18c == out_iindex_1 ? out_prepend_79 : _GEN_3429;
  wire [31:0] _GEN_3431 = 9'h18d == out_iindex_1 ? out_prepend_79 : _GEN_3430;
  wire [31:0] _GEN_3432 = 9'h18e == out_iindex_1 ? out_prepend_79 : _GEN_3431;
  wire [31:0] _GEN_3433 = 9'h18f == out_iindex_1 ? out_prepend_79 : _GEN_3432;
  wire [31:0] _GEN_3434 = 9'h190 == out_iindex_1 ? out_prepend_79 : _GEN_3433;
  wire [31:0] _GEN_3435 = 9'h191 == out_iindex_1 ? out_prepend_79 : _GEN_3434;
  wire [31:0] _GEN_3436 = 9'h192 == out_iindex_1 ? out_prepend_79 : _GEN_3435;
  wire [31:0] _GEN_3437 = 9'h193 == out_iindex_1 ? out_prepend_79 : _GEN_3436;
  wire [31:0] _GEN_3438 = 9'h194 == out_iindex_1 ? out_prepend_79 : _GEN_3437;
  wire [31:0] _GEN_3439 = 9'h195 == out_iindex_1 ? out_prepend_79 : _GEN_3438;
  wire [31:0] _GEN_3440 = 9'h196 == out_iindex_1 ? out_prepend_79 : _GEN_3439;
  wire [31:0] _GEN_3441 = 9'h197 == out_iindex_1 ? out_prepend_79 : _GEN_3440;
  wire [31:0] _GEN_3442 = 9'h198 == out_iindex_1 ? out_prepend_79 : _GEN_3441;
  wire [31:0] _GEN_3443 = 9'h199 == out_iindex_1 ? out_prepend_79 : _GEN_3442;
  wire [31:0] _GEN_3444 = 9'h19a == out_iindex_1 ? out_prepend_79 : _GEN_3443;
  wire [31:0] _GEN_3445 = 9'h19b == out_iindex_1 ? out_prepend_79 : _GEN_3444;
  wire [31:0] _GEN_3446 = 9'h19c == out_iindex_1 ? out_prepend_79 : _GEN_3445;
  wire [31:0] _GEN_3447 = 9'h19d == out_iindex_1 ? out_prepend_79 : _GEN_3446;
  wire [31:0] _GEN_3448 = 9'h19e == out_iindex_1 ? out_prepend_79 : _GEN_3447;
  wire [31:0] _GEN_3449 = 9'h19f == out_iindex_1 ? out_prepend_79 : _GEN_3448;
  wire [31:0] _GEN_3450 = 9'h1a0 == out_iindex_1 ? out_prepend_79 : _GEN_3449;
  wire [31:0] _GEN_3451 = 9'h1a1 == out_iindex_1 ? out_prepend_79 : _GEN_3450;
  wire [31:0] _GEN_3452 = 9'h1a2 == out_iindex_1 ? out_prepend_79 : _GEN_3451;
  wire [31:0] _GEN_3453 = 9'h1a3 == out_iindex_1 ? out_prepend_79 : _GEN_3452;
  wire [31:0] _GEN_3454 = 9'h1a4 == out_iindex_1 ? out_prepend_79 : _GEN_3453;
  wire [31:0] _GEN_3455 = 9'h1a5 == out_iindex_1 ? out_prepend_79 : _GEN_3454;
  wire [31:0] _GEN_3456 = 9'h1a6 == out_iindex_1 ? out_prepend_79 : _GEN_3455;
  wire [31:0] _GEN_3457 = 9'h1a7 == out_iindex_1 ? out_prepend_79 : _GEN_3456;
  wire [31:0] _GEN_3458 = 9'h1a8 == out_iindex_1 ? out_prepend_79 : _GEN_3457;
  wire [31:0] _GEN_3459 = 9'h1a9 == out_iindex_1 ? out_prepend_79 : _GEN_3458;
  wire [31:0] _GEN_3460 = 9'h1aa == out_iindex_1 ? out_prepend_79 : _GEN_3459;
  wire [31:0] _GEN_3461 = 9'h1ab == out_iindex_1 ? out_prepend_79 : _GEN_3460;
  wire [31:0] _GEN_3462 = 9'h1ac == out_iindex_1 ? out_prepend_79 : _GEN_3461;
  wire [31:0] _GEN_3463 = 9'h1ad == out_iindex_1 ? out_prepend_79 : _GEN_3462;
  wire [31:0] _GEN_3464 = 9'h1ae == out_iindex_1 ? out_prepend_79 : _GEN_3463;
  wire [31:0] _GEN_3465 = 9'h1af == out_iindex_1 ? out_prepend_79 : _GEN_3464;
  wire [31:0] _GEN_3466 = 9'h1b0 == out_iindex_1 ? out_prepend_79 : _GEN_3465;
  wire [31:0] _GEN_3467 = 9'h1b1 == out_iindex_1 ? out_prepend_79 : _GEN_3466;
  wire [31:0] _GEN_3468 = 9'h1b2 == out_iindex_1 ? out_prepend_79 : _GEN_3467;
  wire [31:0] _GEN_3469 = 9'h1b3 == out_iindex_1 ? out_prepend_79 : _GEN_3468;
  wire [31:0] _GEN_3470 = 9'h1b4 == out_iindex_1 ? out_prepend_79 : _GEN_3469;
  wire [31:0] _GEN_3471 = 9'h1b5 == out_iindex_1 ? out_prepend_79 : _GEN_3470;
  wire [31:0] _GEN_3472 = 9'h1b6 == out_iindex_1 ? out_prepend_79 : _GEN_3471;
  wire [31:0] _GEN_3473 = 9'h1b7 == out_iindex_1 ? out_prepend_79 : _GEN_3472;
  wire [31:0] _GEN_3474 = 9'h1b8 == out_iindex_1 ? out_prepend_79 : _GEN_3473;
  wire [31:0] _GEN_3475 = 9'h1b9 == out_iindex_1 ? out_prepend_79 : _GEN_3474;
  wire [31:0] _GEN_3476 = 9'h1ba == out_iindex_1 ? out_prepend_79 : _GEN_3475;
  wire [31:0] _GEN_3477 = 9'h1bb == out_iindex_1 ? out_prepend_79 : _GEN_3476;
  wire [31:0] _GEN_3478 = 9'h1bc == out_iindex_1 ? out_prepend_79 : _GEN_3477;
  wire [31:0] _GEN_3479 = 9'h1bd == out_iindex_1 ? out_prepend_79 : _GEN_3478;
  wire [31:0] _GEN_3480 = 9'h1be == out_iindex_1 ? out_prepend_79 : _GEN_3479;
  wire [31:0] _GEN_3481 = 9'h1bf == out_iindex_1 ? out_prepend_79 : _GEN_3480;
  wire [31:0] _GEN_3482 = 9'h1c0 == out_iindex_1 ? out_prepend_79 : _GEN_3481;
  wire [31:0] _GEN_3483 = 9'h1c1 == out_iindex_1 ? out_prepend_79 : _GEN_3482;
  wire [31:0] _GEN_3484 = 9'h1c2 == out_iindex_1 ? out_prepend_79 : _GEN_3483;
  wire [31:0] _GEN_3485 = 9'h1c3 == out_iindex_1 ? out_prepend_79 : _GEN_3484;
  wire [31:0] _GEN_3486 = 9'h1c4 == out_iindex_1 ? out_prepend_79 : _GEN_3485;
  wire [31:0] _GEN_3487 = 9'h1c5 == out_iindex_1 ? out_prepend_79 : _GEN_3486;
  wire [31:0] _GEN_3488 = 9'h1c6 == out_iindex_1 ? out_prepend_79 : _GEN_3487;
  wire [31:0] _GEN_3489 = 9'h1c7 == out_iindex_1 ? out_prepend_79 : _GEN_3488;
  wire [31:0] _GEN_3490 = 9'h1c8 == out_iindex_1 ? out_prepend_79 : _GEN_3489;
  wire [31:0] _GEN_3491 = 9'h1c9 == out_iindex_1 ? out_prepend_79 : _GEN_3490;
  wire [31:0] _GEN_3492 = 9'h1ca == out_iindex_1 ? out_prepend_79 : _GEN_3491;
  wire [31:0] _GEN_3493 = 9'h1cb == out_iindex_1 ? out_prepend_79 : _GEN_3492;
  wire [31:0] _GEN_3494 = 9'h1cc == out_iindex_1 ? out_prepend_79 : _GEN_3493;
  wire [31:0] _GEN_3495 = 9'h1cd == out_iindex_1 ? out_prepend_79 : _GEN_3494;
  wire [31:0] _GEN_3496 = 9'h1ce == out_iindex_1 ? out_prepend_79 : _GEN_3495;
  wire [31:0] _GEN_3497 = 9'h1cf == out_iindex_1 ? out_prepend_79 : _GEN_3496;
  wire [31:0] _GEN_3498 = 9'h1d0 == out_iindex_1 ? out_prepend_79 : _GEN_3497;
  wire [31:0] _GEN_3499 = 9'h1d1 == out_iindex_1 ? out_prepend_79 : _GEN_3498;
  wire [31:0] _GEN_3500 = 9'h1d2 == out_iindex_1 ? out_prepend_79 : _GEN_3499;
  wire [31:0] _GEN_3501 = 9'h1d3 == out_iindex_1 ? out_prepend_79 : _GEN_3500;
  wire [31:0] _GEN_3502 = 9'h1d4 == out_iindex_1 ? out_prepend_79 : _GEN_3501;
  wire [31:0] _GEN_3503 = 9'h1d5 == out_iindex_1 ? out_prepend_79 : _GEN_3502;
  wire [31:0] _GEN_3504 = 9'h1d6 == out_iindex_1 ? out_prepend_79 : _GEN_3503;
  wire [31:0] _GEN_3505 = 9'h1d7 == out_iindex_1 ? out_prepend_79 : _GEN_3504;
  wire [31:0] _GEN_3506 = 9'h1d8 == out_iindex_1 ? out_prepend_79 : _GEN_3505;
  wire [31:0] _GEN_3507 = 9'h1d9 == out_iindex_1 ? out_prepend_79 : _GEN_3506;
  wire [31:0] _GEN_3508 = 9'h1da == out_iindex_1 ? out_prepend_79 : _GEN_3507;
  wire [31:0] _GEN_3509 = 9'h1db == out_iindex_1 ? out_prepend_79 : _GEN_3508;
  wire [31:0] _GEN_3510 = 9'h1dc == out_iindex_1 ? out_prepend_79 : _GEN_3509;
  wire [31:0] _GEN_3511 = 9'h1dd == out_iindex_1 ? out_prepend_79 : _GEN_3510;
  wire [31:0] _GEN_3512 = 9'h1de == out_iindex_1 ? out_prepend_79 : _GEN_3511;
  wire [31:0] _GEN_3513 = 9'h1df == out_iindex_1 ? out_prepend_79 : _GEN_3512;
  wire [31:0] _GEN_3514 = 9'h1e0 == out_iindex_1 ? out_prepend_79 : _GEN_3513;
  wire [31:0] _GEN_3515 = 9'h1e1 == out_iindex_1 ? out_prepend_79 : _GEN_3514;
  wire [31:0] _GEN_3516 = 9'h1e2 == out_iindex_1 ? out_prepend_79 : _GEN_3515;
  wire [31:0] _GEN_3517 = 9'h1e3 == out_iindex_1 ? out_prepend_79 : _GEN_3516;
  wire [31:0] _GEN_3518 = 9'h1e4 == out_iindex_1 ? out_prepend_79 : _GEN_3517;
  wire [31:0] _GEN_3519 = 9'h1e5 == out_iindex_1 ? out_prepend_79 : _GEN_3518;
  wire [31:0] _GEN_3520 = 9'h1e6 == out_iindex_1 ? out_prepend_79 : _GEN_3519;
  wire [31:0] _GEN_3521 = 9'h1e7 == out_iindex_1 ? out_prepend_79 : _GEN_3520;
  wire [31:0] _GEN_3522 = 9'h1e8 == out_iindex_1 ? out_prepend_79 : _GEN_3521;
  wire [31:0] _GEN_3523 = 9'h1e9 == out_iindex_1 ? out_prepend_79 : _GEN_3522;
  wire [31:0] _GEN_3524 = 9'h1ea == out_iindex_1 ? out_prepend_79 : _GEN_3523;
  wire [31:0] _GEN_3525 = 9'h1eb == out_iindex_1 ? out_prepend_79 : _GEN_3524;
  wire [31:0] _GEN_3526 = 9'h1ec == out_iindex_1 ? out_prepend_79 : _GEN_3525;
  wire [31:0] _GEN_3527 = 9'h1ed == out_iindex_1 ? out_prepend_79 : _GEN_3526;
  wire [31:0] _GEN_3528 = 9'h1ee == out_iindex_1 ? out_prepend_79 : _GEN_3527;
  wire [31:0] _GEN_3529 = 9'h1ef == out_iindex_1 ? out_prepend_79 : _GEN_3528;
  wire [31:0] _GEN_3530 = 9'h1f0 == out_iindex_1 ? out_prepend_79 : _GEN_3529;
  wire [31:0] _GEN_3531 = 9'h1f1 == out_iindex_1 ? out_prepend_79 : _GEN_3530;
  wire [31:0] _GEN_3532 = 9'h1f2 == out_iindex_1 ? out_prepend_79 : _GEN_3531;
  wire [31:0] _GEN_3533 = 9'h1f3 == out_iindex_1 ? out_prepend_79 : _GEN_3532;
  wire [31:0] _GEN_3534 = 9'h1f4 == out_iindex_1 ? out_prepend_79 : _GEN_3533;
  wire [31:0] _GEN_3535 = 9'h1f5 == out_iindex_1 ? out_prepend_79 : _GEN_3534;
  wire [31:0] _GEN_3536 = 9'h1f6 == out_iindex_1 ? out_prepend_79 : _GEN_3535;
  wire [31:0] _GEN_3537 = 9'h1f7 == out_iindex_1 ? out_prepend_79 : _GEN_3536;
  wire [31:0] _GEN_3538 = 9'h1f8 == out_iindex_1 ? out_prepend_79 : _GEN_3537;
  wire [31:0] _GEN_3539 = 9'h1f9 == out_iindex_1 ? out_prepend_79 : _GEN_3538;
  wire [31:0] _GEN_3540 = 9'h1fa == out_iindex_1 ? out_prepend_79 : _GEN_3539;
  wire [31:0] _GEN_3541 = 9'h1fb == out_iindex_1 ? out_prepend_79 : _GEN_3540;
  wire [31:0] _GEN_3542 = 9'h1fc == out_iindex_1 ? out_prepend_79 : _GEN_3541;
  wire [31:0] _GEN_3543 = 9'h1fd == out_iindex_1 ? out_prepend_79 : _GEN_3542;
  wire [31:0] _GEN_3544 = 9'h1fe == out_iindex_1 ? out_prepend_79 : _GEN_3543;
  wire [31:0] _GEN_3545 = 9'h1ff == out_iindex_1 ? out_prepend_79 : _GEN_3544;
  wire [1:0] _GEN_3627 = commandRegBadHaltResume ? 2'h0 : 2'h2;
  wire [1:0] _GEN_3633 = ~goReg & out_f_woready_647 ? 2'h0 : ctrlStateReg;
  wire [1:0] _GEN_3634 = out_f_woready_941 ? 2'h0 : _GEN_3633;
  wire  _T_1393 = ctrlStateReg == 2'h3;
  wire  _GEN_3894 = _errorBusy_T & ~_T_1383;
  
  
  AsyncResetSynchronizerShiftReg_w1_d3_i0 hartIsInResetSync_0_debug_hartReset_0 (
    .clock(hartIsInResetSync_0_debug_hartReset_0_clock),
    .reset(hartIsInResetSync_0_debug_hartReset_0_reset),
    .io_d(hartIsInResetSync_0_debug_hartReset_0_io_d),
    .io_q(hartIsInResetSync_0_debug_hartReset_0_io_q)
  );
  assign auto_tl_in_a_ready = auto_tl_in_d_ready;
  assign auto_tl_in_d_valid = auto_tl_in_a_valid;
  assign auto_tl_in_d_bits_opcode = {{2'd0}, in_1_bits_read};
  assign auto_tl_in_d_bits_size = auto_tl_in_a_bits_size;
  assign auto_tl_in_d_bits_source = auto_tl_in_a_bits_source;
  assign auto_tl_in_d_bits_data = _GEN_3033 ? _GEN_3545 : 32'h0;
  assign auto_dmi_in_a_ready = auto_dmi_in_d_ready;
  assign auto_dmi_in_d_valid = auto_dmi_in_a_valid;
  assign auto_dmi_in_d_bits_opcode = {{2'd0}, in_bits_read};
  assign auto_dmi_in_d_bits_size = auto_dmi_in_a_bits_size;
  assign auto_dmi_in_d_bits_source = auto_dmi_in_a_bits_source;
  assign auto_dmi_in_d_bits_data = _GEN_296 ? _GEN_328 : 32'h0;
  assign io_innerCtrl_ready = 1'h1;
  assign io_hgDebugInt_0 = hrDebugIntReg_0;
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = auto_dmi_in_d_ready;
  assign monitor_io_in_a_valid = auto_dmi_in_a_valid;
  assign monitor_io_in_a_bits_opcode = auto_dmi_in_a_bits_opcode;
  assign monitor_io_in_a_bits_param = auto_dmi_in_a_bits_param;
  assign monitor_io_in_a_bits_size = auto_dmi_in_a_bits_size;
  assign monitor_io_in_a_bits_source = auto_dmi_in_a_bits_source;
  assign monitor_io_in_a_bits_address = auto_dmi_in_a_bits_address;
  assign monitor_io_in_a_bits_mask = auto_dmi_in_a_bits_mask;
  assign monitor_io_in_a_bits_corrupt = auto_dmi_in_a_bits_corrupt;
  assign monitor_io_in_d_ready = auto_dmi_in_d_ready;
  assign monitor_io_in_d_valid = auto_dmi_in_a_valid;
  assign monitor_io_in_d_bits_opcode = {{2'd0}, in_bits_read};
  assign monitor_io_in_d_bits_size = auto_dmi_in_a_bits_size;
  assign monitor_io_in_d_bits_source = auto_dmi_in_a_bits_source;
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_a_ready = auto_tl_in_d_ready;
  assign monitor_1_io_in_a_valid = auto_tl_in_a_valid;
  assign monitor_1_io_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
  assign monitor_1_io_in_a_bits_param = auto_tl_in_a_bits_param;
  assign monitor_1_io_in_a_bits_size = auto_tl_in_a_bits_size;
  assign monitor_1_io_in_a_bits_source = auto_tl_in_a_bits_source;
  assign monitor_1_io_in_a_bits_address = auto_tl_in_a_bits_address;
  assign monitor_1_io_in_a_bits_mask = auto_tl_in_a_bits_mask;
  assign monitor_1_io_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
  assign monitor_1_io_in_d_ready = auto_tl_in_d_ready;
  assign monitor_1_io_in_d_valid = auto_tl_in_a_valid;
  assign monitor_1_io_in_d_bits_opcode = {{2'd0}, in_1_bits_read};
  assign monitor_1_io_in_d_bits_size = auto_tl_in_a_bits_size;
  assign monitor_1_io_in_d_bits_source = auto_tl_in_a_bits_source;
  assign hartIsInResetSync_0_debug_hartReset_0_clock = clock;
  assign hartIsInResetSync_0_debug_hartReset_0_reset = reset;
  assign hartIsInResetSync_0_debug_hartReset_0_io_d = io_hartIsInReset_0;
  always @(posedge clock) begin
    haltedBitRegs <= _GEN_65[0];
    resumeReqRegs <= _GEN_66[0];
    if (_T_1) begin
      haveResetBitRegs <= 1'h0;
    end else if (_T_4 & io_innerCtrl_bits_ackhavereset) begin
      haveResetBitRegs <= haveResetBitRegs & _resumeAcks_T_1 | hartIsInResetSync_0;
    end else begin
      haveResetBitRegs <= haveResetBitRegs | hartIsInResetSync_0;
    end
    if (reset) begin
      hrmaskReg_0 <= 1'h0;
    end else if (~io_dmactive) begin
      hrmaskReg_0 <= 1'h0;
    end else if (_T_4) begin
      hrmaskReg_0 <= io_innerCtrl_bits_hrmask_0;
    end
    if (_T_1) begin
      ABSTRACTCSReg_cmderr <= 3'h0;
    end else if (errorBusy) begin
      ABSTRACTCSReg_cmderr <= 3'h1;
    end else if (errorException) begin
      ABSTRACTCSReg_cmderr <= 3'h3;
    end else if (errorUnsupported) begin
      ABSTRACTCSReg_cmderr <= 3'h2;
    end else begin
      ABSTRACTCSReg_cmderr <= _GEN_38;
    end
    if (_T_1) begin
      ctrlStateReg <= 2'h0;
    end else if (ABSTRACTCSWrEnLegal) begin
      if (wrAccessRegisterCommand | regAccessRegisterCommand) begin
        ctrlStateReg <= 2'h1;
      end
    end else if (ctrlStateReg == 2'h1) begin
      if (commandRegIsUnsupported) begin
        ctrlStateReg <= 2'h0;
      end else begin
        ctrlStateReg <= _GEN_3627;
      end
    end else if (ctrlStateReg == 2'h2) begin
      ctrlStateReg <= _GEN_3634;
    end
    if (_T_1) begin
      COMMANDRdData_cmdtype <= 8'h0;
    end else if (COMMANDWrEn) begin
      COMMANDRdData_cmdtype <= COMMANDWrData_cmdtype;
    end
    if (_T_1) begin
      COMMANDRdData_control <= 24'h0;
    end else if (COMMANDWrEn) begin
      COMMANDRdData_control <= COMMANDWrData_control;
    end
    if (_T_1) begin
      ABSTRACTAUTOReg_autoexecdata <= 12'h0;
    end else if (out_f_woready_4 & ABSTRACTCSWrEnLegal) begin
      ABSTRACTAUTOReg_autoexecdata <= _ABSTRACTAUTOReg_autoexecdata_T;
    end
    if (_T_1) begin
      ABSTRACTAUTOReg_autoexecprogbuf <= 16'h0;
    end else if (out_f_woready_6 & ABSTRACTCSWrEnLegal) begin
      ABSTRACTAUTOReg_autoexecprogbuf <= ABSTRACTAUTOWrData_autoexecprogbuf;
    end
    if (_T_1) begin
      abstractDataMem_0 <= 8'h0;
    end else if (out_f_wivalid_503) begin
      abstractDataMem_0 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_92 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_92) begin
        abstractDataMem_0 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      abstractDataMem_1 <= 8'h0;
    end else if (out_f_wivalid_504) begin
      abstractDataMem_1 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_93 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_93) begin
        abstractDataMem_1 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      abstractDataMem_2 <= 8'h0;
    end else if (out_f_wivalid_505) begin
      abstractDataMem_2 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_94 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_94) begin
        abstractDataMem_2 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      abstractDataMem_3 <= 8'h0;
    end else if (out_f_wivalid_506) begin
      abstractDataMem_3 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_95 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_95) begin
        abstractDataMem_3 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_0 <= 8'h0;
    end else if (out_f_wivalid_768) begin
      programBufferMem_0 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_27 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_27) begin
        programBufferMem_0 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_1 <= 8'h0;
    end else if (out_f_wivalid_769) begin
      programBufferMem_1 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_28 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_28) begin
        programBufferMem_1 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_2 <= 8'h0;
    end else if (out_f_wivalid_770) begin
      programBufferMem_2 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_29 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_29) begin
        programBufferMem_2 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_3 <= 8'h0;
    end else if (out_f_wivalid_771) begin
      programBufferMem_3 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_30 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_30) begin
        programBufferMem_3 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_4 <= 8'h0;
    end else if (out_f_wivalid_885) begin
      programBufferMem_4 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_19 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_19) begin
        programBufferMem_4 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_5 <= 8'h0;
    end else if (out_f_wivalid_886) begin
      programBufferMem_5 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_20 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_20) begin
        programBufferMem_5 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_6 <= 8'h0;
    end else if (out_f_wivalid_887) begin
      programBufferMem_6 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_21 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_21) begin
        programBufferMem_6 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_7 <= 8'h0;
    end else if (out_f_wivalid_888) begin
      programBufferMem_7 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_22 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_22) begin
        programBufferMem_7 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_8 <= 8'h0;
    end else if (out_f_wivalid_1143) begin
      programBufferMem_8 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_31 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_31) begin
        programBufferMem_8 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_9 <= 8'h0;
    end else if (out_f_wivalid_1144) begin
      programBufferMem_9 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_32 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_32) begin
        programBufferMem_9 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_10 <= 8'h0;
    end else if (out_f_wivalid_1145) begin
      programBufferMem_10 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_33 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_33) begin
        programBufferMem_10 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_11 <= 8'h0;
    end else if (out_f_wivalid_1146) begin
      programBufferMem_11 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_34 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_34) begin
        programBufferMem_11 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_12 <= 8'h0;
    end else if (out_f_wivalid_300) begin
      programBufferMem_12 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_74 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_74) begin
        programBufferMem_12 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_13 <= 8'h0;
    end else if (out_f_wivalid_301) begin
      programBufferMem_13 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_75 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_75) begin
        programBufferMem_13 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_14 <= 8'h0;
    end else if (out_f_wivalid_302) begin
      programBufferMem_14 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_76 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_76) begin
        programBufferMem_14 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_15 <= 8'h0;
    end else if (out_f_wivalid_303) begin
      programBufferMem_15 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_77 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_77) begin
        programBufferMem_15 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_16 <= 8'h0;
    end else if (out_f_wivalid_567) begin
      programBufferMem_16 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_87 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_87) begin
        programBufferMem_16 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_17 <= 8'h0;
    end else if (out_f_wivalid_568) begin
      programBufferMem_17 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_88 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_88) begin
        programBufferMem_17 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_18 <= 8'h0;
    end else if (out_f_wivalid_569) begin
      programBufferMem_18 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_89 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_89) begin
        programBufferMem_18 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_19 <= 8'h0;
    end else if (out_f_wivalid_570) begin
      programBufferMem_19 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_90 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_90) begin
        programBufferMem_19 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_20 <= 8'h0;
    end else if (out_f_wivalid_796) begin
      programBufferMem_20 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_7 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_7) begin
        programBufferMem_20 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_21 <= 8'h0;
    end else if (out_f_wivalid_797) begin
      programBufferMem_21 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_8 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_8) begin
        programBufferMem_21 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_22 <= 8'h0;
    end else if (out_f_wivalid_798) begin
      programBufferMem_22 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_9 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_9) begin
        programBufferMem_22 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_23 <= 8'h0;
    end else if (out_f_wivalid_799) begin
      programBufferMem_23 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_10 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_10) begin
        programBufferMem_23 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_24 <= 8'h0;
    end else if (out_f_wivalid_1091) begin
      programBufferMem_24 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_15 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_15) begin
        programBufferMem_24 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_25 <= 8'h0;
    end else if (out_f_wivalid_1092) begin
      programBufferMem_25 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_16 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_16) begin
        programBufferMem_25 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_26 <= 8'h0;
    end else if (out_f_wivalid_1093) begin
      programBufferMem_26 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_17 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_17) begin
        programBufferMem_26 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_27 <= 8'h0;
    end else if (out_f_wivalid_1094) begin
      programBufferMem_27 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_18 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_18) begin
        programBufferMem_27 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_28 <= 8'h0;
    end else if (out_f_wivalid_1259) begin
      programBufferMem_28 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_70 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_70) begin
        programBufferMem_28 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_29 <= 8'h0;
    end else if (out_f_wivalid_1260) begin
      programBufferMem_29 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_71 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_71) begin
        programBufferMem_29 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_30 <= 8'h0;
    end else if (out_f_wivalid_1261) begin
      programBufferMem_30 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_72 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_72) begin
        programBufferMem_30 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_31 <= 8'h0;
    end else if (out_f_wivalid_1262) begin
      programBufferMem_31 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_73 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_73) begin
        programBufferMem_31 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_32 <= 8'h0;
    end else if (out_f_wivalid_276) begin
      programBufferMem_32 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_82 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_82) begin
        programBufferMem_32 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_33 <= 8'h0;
    end else if (out_f_wivalid_277) begin
      programBufferMem_33 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_83 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_83) begin
        programBufferMem_33 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_34 <= 8'h0;
    end else if (out_f_wivalid_278) begin
      programBufferMem_34 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_84 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_84) begin
        programBufferMem_34 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_35 <= 8'h0;
    end else if (out_f_wivalid_279) begin
      programBufferMem_35 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_85 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_85) begin
        programBufferMem_35 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_36 <= 8'h0;
    end else if (out_f_wivalid_140) begin
      programBufferMem_36 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_23 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_23) begin
        programBufferMem_36 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_37 <= 8'h0;
    end else if (out_f_wivalid_141) begin
      programBufferMem_37 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_24 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_24) begin
        programBufferMem_37 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_38 <= 8'h0;
    end else if (out_f_wivalid_142) begin
      programBufferMem_38 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_25 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_25) begin
        programBufferMem_38 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_39 <= 8'h0;
    end else if (out_f_wivalid_143) begin
      programBufferMem_39 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_26 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_26) begin
        programBufferMem_39 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_40 <= 8'h0;
    end else if (out_f_wivalid_1018) begin
      programBufferMem_40 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready) begin
        programBufferMem_40 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_41 <= 8'h0;
    end else if (out_f_wivalid_1019) begin
      programBufferMem_41 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_1 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_1) begin
        programBufferMem_41 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_42 <= 8'h0;
    end else if (out_f_wivalid_1020) begin
      programBufferMem_42 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_2 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_2) begin
        programBufferMem_42 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_43 <= 8'h0;
    end else if (out_f_wivalid_1021) begin
      programBufferMem_43 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_3 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_3) begin
        programBufferMem_43 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_44 <= 8'h0;
    end else if (out_f_wivalid_724) begin
      programBufferMem_44 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_78 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_78) begin
        programBufferMem_44 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_45 <= 8'h0;
    end else if (out_f_wivalid_725) begin
      programBufferMem_45 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_79 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_79) begin
        programBufferMem_45 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_46 <= 8'h0;
    end else if (out_f_wivalid_726) begin
      programBufferMem_46 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_80 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_80) begin
        programBufferMem_46 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_47 <= 8'h0;
    end else if (out_f_wivalid_727) begin
      programBufferMem_47 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_81 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_81) begin
        programBufferMem_47 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_48 <= 8'h0;
    end else if (out_f_wivalid_409) begin
      programBufferMem_48 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_66 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_66) begin
        programBufferMem_48 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_49 <= 8'h0;
    end else if (out_f_wivalid_410) begin
      programBufferMem_49 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_67 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_67) begin
        programBufferMem_49 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_50 <= 8'h0;
    end else if (out_f_wivalid_411) begin
      programBufferMem_50 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_68 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_68) begin
        programBufferMem_50 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_51 <= 8'h0;
    end else if (out_f_wivalid_412) begin
      programBufferMem_51 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_69 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_69) begin
        programBufferMem_51 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_52 <= 8'h0;
    end else if (out_f_wivalid_332) begin
      programBufferMem_52 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_35 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_35) begin
        programBufferMem_52 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_53 <= 8'h0;
    end else if (out_f_wivalid_333) begin
      programBufferMem_53 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_36 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_36) begin
        programBufferMem_53 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_54 <= 8'h0;
    end else if (out_f_wivalid_334) begin
      programBufferMem_54 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_37 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_37) begin
        programBufferMem_54 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_55 <= 8'h0;
    end else if (out_f_wivalid_335) begin
      programBufferMem_55 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_38 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_38) begin
        programBufferMem_55 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_56 <= 8'h0;
    end else if (out_f_wivalid_1267) begin
      programBufferMem_56 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_11 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_11) begin
        programBufferMem_56 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_57 <= 8'h0;
    end else if (out_f_wivalid_1268) begin
      programBufferMem_57 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_12 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_12) begin
        programBufferMem_57 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_58 <= 8'h0;
    end else if (out_f_wivalid_1269) begin
      programBufferMem_58 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_13 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_13) begin
        programBufferMem_58 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_59 <= 8'h0;
    end else if (out_f_wivalid_1270) begin
      programBufferMem_59 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_14 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_14) begin
        programBufferMem_59 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      programBufferMem_60 <= 8'h0;
    end else if (out_f_wivalid_833) begin
      programBufferMem_60 <= auto_tl_in_a_bits_data[7:0];
    end else if (out_f_woready_96 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_96) begin
        programBufferMem_60 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_1) begin
      programBufferMem_61 <= 8'h0;
    end else if (out_f_wivalid_834) begin
      programBufferMem_61 <= auto_tl_in_a_bits_data[15:8];
    end else if (out_f_woready_97 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_97) begin
        programBufferMem_61 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_1) begin
      programBufferMem_62 <= 8'h0;
    end else if (out_f_wivalid_835) begin
      programBufferMem_62 <= auto_tl_in_a_bits_data[23:16];
    end else if (out_f_woready_98 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_98) begin
        programBufferMem_62 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_1) begin
      programBufferMem_63 <= 8'h0;
    end else if (out_f_wivalid_836) begin
      programBufferMem_63 <= auto_tl_in_a_bits_data[31:24];
    end else if (out_f_woready_99 & ABSTRACTCSWrEnLegal) begin
      if (out_f_woready_99) begin
        programBufferMem_63 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_1) begin
      goReg <= 1'h0;
    end else begin
      goReg <= _GEN_398;
    end
    if (goAbstract) begin
      if (accessRegisterCommandReg_transfer) begin
        if (accessRegisterCommandReg_write) begin
          abstractGeneratedMem_0 <= _abstractGeneratedMem_0_T;
        end else begin
          abstractGeneratedMem_0 <= _abstractGeneratedMem_0_T_1;
        end
      end else begin
        abstractGeneratedMem_0 <= 32'h13;
      end
    end
    if (goAbstract) begin
      if (accessRegisterCommandReg_postexec) begin
        abstractGeneratedMem_1 <= 32'h13;
      end else begin
        abstractGeneratedMem_1 <= 32'h100073;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(hartGoingId == 10'h0) & (~_T_1 & ~goAbstract & out_f_woready_470 & ~reset)) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1 & ~goAbstract & out_f_woready_470 & ~reset & ~(hartGoingId == 10'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Unexpected 'GOING' hart.\n    at Debug.scala:1390 assert(hartGoingId === 0.U, \"Unexpected 'GOING' hart.\")//Chisel3 #540 %%x, expected %%x\", hartGoingId, 0.U)\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_342 & (_errorBusy_T & ~_T_1383 & _T_1384 & out_f_woready_941 & _T_341)) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_errorBusy_T & ~_T_1383 & _T_1384 & out_f_woready_941 & _T_341 & _T_342) begin
          $fwrite(32'h80000002,
            "Assertion failed: Unexpected 'EXCEPTION' hart\n    at Debug.scala:1710 assert(hartExceptionId === 0.U, \"Unexpected 'EXCEPTION' hart\")//Chisel3 #540, %%x, expected %%x\", hartExceptionId, 0.U)\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_3894 & ~_T_1384 & _T_1393 & _T_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_3894 & ~_T_1384 & _T_1393 & _T_341) begin
          $fwrite(32'h80000002,
            "Assertion failed: Should not be in custom state unless we need it.\n    at Debug.scala:1715 assert(needCustom.B, \"Should not be in custom state unless we need it.\")\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1 | ~out_f_woready_941 | _T_1384) & _T_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_341 & ~(_T_1 | ~out_f_woready_941 | _T_1384)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Unexpected EXCEPTION write: should only get it in Debug Module EXEC state\n    at Debug.scala:1728 assert ((!io.dmactive || !hartExceptionWrEn || ctrlStateReg === CtrlState(Exec)),\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      hrDebugIntReg_0 <= 1'h0;
    end else if (_T_1) begin
      hrDebugIntReg_0 <= 1'h0;
    end else begin
      hrDebugIntReg_0 <= _T_13;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  haltedBitRegs = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resumeReqRegs = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  haveResetBitRegs = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  hrmaskReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  hrDebugIntReg_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ABSTRACTCSReg_cmderr = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  ctrlStateReg = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  COMMANDRdData_cmdtype = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  COMMANDRdData_control = _RAND_8[23:0];
  _RAND_9 = {1{`RANDOM}};
  ABSTRACTAUTOReg_autoexecdata = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  ABSTRACTAUTOReg_autoexecprogbuf = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  abstractDataMem_0 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  abstractDataMem_1 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  abstractDataMem_2 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  abstractDataMem_3 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  programBufferMem_0 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  programBufferMem_1 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  programBufferMem_2 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  programBufferMem_3 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  programBufferMem_4 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  programBufferMem_5 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  programBufferMem_6 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  programBufferMem_7 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  programBufferMem_8 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  programBufferMem_9 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  programBufferMem_10 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  programBufferMem_11 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  programBufferMem_12 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  programBufferMem_13 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  programBufferMem_14 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  programBufferMem_15 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  programBufferMem_16 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  programBufferMem_17 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  programBufferMem_18 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  programBufferMem_19 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  programBufferMem_20 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  programBufferMem_21 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  programBufferMem_22 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  programBufferMem_23 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  programBufferMem_24 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  programBufferMem_25 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  programBufferMem_26 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  programBufferMem_27 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  programBufferMem_28 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  programBufferMem_29 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  programBufferMem_30 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  programBufferMem_31 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  programBufferMem_32 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  programBufferMem_33 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  programBufferMem_34 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  programBufferMem_35 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  programBufferMem_36 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  programBufferMem_37 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  programBufferMem_38 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  programBufferMem_39 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  programBufferMem_40 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  programBufferMem_41 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  programBufferMem_42 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  programBufferMem_43 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  programBufferMem_44 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  programBufferMem_45 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  programBufferMem_46 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  programBufferMem_47 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  programBufferMem_48 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  programBufferMem_49 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  programBufferMem_50 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  programBufferMem_51 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  programBufferMem_52 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  programBufferMem_53 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  programBufferMem_54 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  programBufferMem_55 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  programBufferMem_56 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  programBufferMem_57 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  programBufferMem_58 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  programBufferMem_59 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  programBufferMem_60 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  programBufferMem_61 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  programBufferMem_62 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  programBufferMem_63 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  goReg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  abstractGeneratedMem_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  abstractGeneratedMem_1 = _RAND_81[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    hrDebugIntReg_0 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule