// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-08-13
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_313
`define RVX_GDEF_313

`define RVX_GDEF_100 None
`define RVX_GDEF_337 8
`define RVX_GDEF_189 3
`define RVX_GDEF_261 0

`define RVX_GDEF_214 5
`define RVX_GDEF_175 0
`define RVX_GDEF_222 0
`define RVX_GDEF_345 16
`define RVX_GDEF_400 20
`define RVX_GDEF_202 21
`define RVX_GDEF_182 22
`define RVX_GDEF_423 23
`define RVX_GDEF_376 24
`define RVX_GDEF_239 28

`define RVX_GDEF_272 5
`define RVX_GDEF_181 0
`define RVX_GDEF_039 16
`define RVX_GDEF_110 4
`define RVX_GDEF_034 1
`define RVX_GDEF_119 1
`define RVX_GDEF_167 1
`define RVX_GDEF_021 1
`define RVX_GDEF_076 1
`define RVX_GDEF_094 3

`endif